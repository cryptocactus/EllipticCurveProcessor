
//256-b_notit Carry Look Ahead Adder with overflow b_notit
//Created b_noty: Colter Sisler, Scott Everitt, Steven Dougherty
//Team: Nighthawk
//Rev: 3.0
//2-22-2017


module sub_256 (
  input [255:0] a,
  input [255:0] b,
  output reg [255:0] sum,
  output wire carry_out_overflow_not
);

wire carry_in_n;
wire signed [255:0] b_not;
reg signed [255:0] g,p;
reg signed [255:0] carry_in;
reg signed [255:1] carry_out;
reg carry_out_overflow;

assign carry_out_overflow_not = ~carry_out_overflow;

assign carry_in_n = 1'b1;

assign b_not = ~b;

always @* begin




carry_out[1] = (((a[0]^b_not[0])&carry_in_n)|(a[0]&b_not[0]));
g[0] = a[0]&b_not[0];
p[0] = a[0]^b_not[0];
sum[0] = p[0]^carry_in_n;
carry_in[0] = carry_in_n;
carry_in[1] = (g[0] | carry_in[0]&p[0]);

g[1] = a[1]&b_not[1];
p[1] = a[1]^b_not[1];
sum[1]= (p[1]^carry_in[1]);
carry_in[2] = (g[1]|carry_in[1]&p[1]);
carry_out[2] = (g[1] | p[1] &(g[0] | carry_in[0]&p[0]));

g[2] = a[2]&b_not[2];
p[2] = a[2]^b_not[2];
sum[2]= (p[2]^carry_in[2]);
carry_in[3] = (g[2]|carry_in[2]&p[2]);
carry_out[3] = (g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])));

g[3] = a[3]&b_not[3];
p[3] = a[3]^b_not[3];
sum[3]= (p[3]^carry_in[3]);
carry_in[4] = (g[3]|carry_in[3]&p[3]);
carry_out[4] = (g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))));
g[4] = a[4]&b_not[4];
p[4] = a[4]^b_not[4];

sum[4]= (p[4]^carry_in[4]);
carry_in[5] = (g[4]|carry_in[4]&p[4]);
carry_out[5] = (g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))));
g[5] = a[5]&b_not[5];
p[5] = a[5]^b_not[5];

sum[5]= (p[5]^carry_in[5]);
carry_in[6] = (g[5]|carry_in[5]&p[5]);
carry_out[6] = (g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))));
g[6] = a[6]&b_not[6];
p[6] = a[6]^b_not[6];

sum[6]= (p[6]^carry_in[6]);
carry_in[7] = (g[6]|carry_in[6]&p[6]);
carry_out[7] = (g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))));
g[7] = a[7]&b_not[7];
p[7] = a[7]^b_not[7];

sum[7]= (p[7]^carry_in[7]);
carry_in[8] = (g[7]|carry_in[7]&p[7]);
carry_out[8] = (g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))));
g[8] = a[8]&b_not[8];
p[8] = a[8]^b_not[8];

sum[8]= (p[8]^carry_in[8]);
carry_in[9] = (g[8]|carry_in[8]&p[8]);
carry_out[9] = (g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))));
g[9] = a[9]&b_not[9];
p[9] = a[9]^b_not[9];

sum[9]= (p[9]^carry_in[9]);
carry_in[10] = (g[9]|carry_in[9]&p[9]);
carry_out[10] = (g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))));
g[10] = a[10]&b_not[10];
p[10] = a[10]^b_not[10];

sum[10]= (p[10]^carry_in[10]);
carry_in[11] = (g[10]|carry_in[10]&p[10]);
carry_out[11] = (g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))));
g[11] = a[11]&b_not[11];
p[11] = a[11]^b_not[11];

sum[11]= (p[11]^carry_in[11]);
carry_in[12] = (g[11]|carry_in[11]&p[11]);
carry_out[12] = (g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))));
g[12] = a[12]&b_not[12];
p[12] = a[12]^b_not[12];

sum[12]= (p[12]^carry_in[12]);
carry_in[13] = (g[12]|carry_in[12]&p[12]);
carry_out[13] = (g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))));
g[13] = a[13]&b_not[13];
p[13] = a[13]^b_not[13];

sum[13]= (p[13]^carry_in[13]);
carry_in[14] = (g[13]|carry_in[13]&p[13]);
carry_out[14] = (g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))));
g[14] = a[14]&b_not[14];
p[14] = a[14]^b_not[14];

sum[14]= (p[14]^carry_in[14]);
carry_in[15] = (g[14]|carry_in[14]&p[14]);
carry_out[15] = (g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))));
g[15] = a[15]&b_not[15];
p[15] = a[15]^b_not[15];

sum[15]= (p[15]^carry_in[15]);
carry_in[16] = (g[15]|carry_in[15]&p[15]);
carry_out[16] = (g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))));
g[16] = a[16]&b_not[16];
p[16] = a[16]^b_not[16];

sum[16]= (p[16]^carry_in[16]);
carry_in[17] = (g[16]|carry_in[16]&p[16]);
carry_out[17] = (g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))));
g[17] = a[17]&b_not[17];
p[17] = a[17]^b_not[17];

sum[17]= (p[17]^carry_in[17]);
carry_in[18] = (g[17]|carry_in[17]&p[17]);
carry_out[18] = (g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))));
g[18] = a[18]&b_not[18];
p[18] = a[18]^b_not[18];

sum[18]= (p[18]^carry_in[18]);
carry_in[19] = (g[18]|carry_in[18]&p[18]);
carry_out[19] = (g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))));
g[19] = a[19]&b_not[19];
p[19] = a[19]^b_not[19];

sum[19]= (p[19]^carry_in[19]);
carry_in[20] = (g[19]|carry_in[19]&p[19]);
carry_out[20] = (g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))));
g[20] = a[20]&b_not[20];
p[20] = a[20]^b_not[20];

sum[20]= (p[20]^carry_in[20]);
carry_in[21] = (g[20]|carry_in[20]&p[20]);
carry_out[21] = (g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))));
g[21] = a[21]&b_not[21];
p[21] = a[21]^b_not[21];

sum[21]= (p[21]^carry_in[21]);
carry_in[22] = (g[21]|carry_in[21]&p[21]);
carry_out[22] = (g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))));
g[22] = a[22]&b_not[22];
p[22] = a[22]^b_not[22];

sum[22]= (p[22]^carry_in[22]);
carry_in[23] = (g[22]|carry_in[22]&p[22]);
carry_out[23] = (g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))));
g[23] = a[23]&b_not[23];
p[23] = a[23]^b_not[23];

sum[23]= (p[23]^carry_in[23]);
carry_in[24] = (g[23]|carry_in[23]&p[23]);
carry_out[24] = (g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))));
g[24] = a[24]&b_not[24];
p[24] = a[24]^b_not[24];

sum[24]= (p[24]^carry_in[24]);
carry_in[25] = (g[24]|carry_in[24]&p[24]);
carry_out[25] = (g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))));
g[25] = a[25]&b_not[25];
p[25] = a[25]^b_not[25];

sum[25]= (p[25]^carry_in[25]);
carry_in[26] = (g[25]|carry_in[25]&p[25]);
carry_out[26] = (g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))));
g[26] = a[26]&b_not[26];
p[26] = a[26]^b_not[26];

sum[26]= (p[26]^carry_in[26]);
carry_in[27] = (g[26]|carry_in[26]&p[26]);
carry_out[27] = (g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))));
g[27] = a[27]&b_not[27];
p[27] = a[27]^b_not[27];

sum[27]= (p[27]^carry_in[27]);
carry_in[28] = (g[27]|carry_in[27]&p[27]);
carry_out[28] = (g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))));
g[28] = a[28]&b_not[28];
p[28] = a[28]^b_not[28];

sum[28]= (p[28]^carry_in[28]);
carry_in[29] = (g[28]|carry_in[28]&p[28]);
carry_out[29] = (g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))));
g[29] = a[29]&b_not[29];
p[29] = a[29]^b_not[29];

sum[29]= (p[29]^carry_in[29]);
carry_in[30] = (g[29]|carry_in[29]&p[29]);
carry_out[30] = (g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))));
g[30] = a[30]&b_not[30];
p[30] = a[30]^b_not[30];

sum[30]= (p[30]^carry_in[30]);
carry_in[31] = (g[30]|carry_in[30]&p[30]);
carry_out[31] = (g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))));
g[31] = a[31]&b_not[31];
p[31] = a[31]^b_not[31];

sum[31]= (p[31]^carry_in[31]);
carry_in[32] = (g[31]|carry_in[31]&p[31]);
carry_out[32] = (g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))));
g[32] = a[32]&b_not[32];
p[32] = a[32]^b_not[32];

sum[32]= (p[32]^carry_in[32]);
carry_in[33] = (g[32]|carry_in[32]&p[32]);
carry_out[33] = (g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))));
g[33] = a[33]&b_not[33];
p[33] = a[33]^b_not[33];

sum[33]= (p[33]^carry_in[33]);
carry_in[34] = (g[33]|carry_in[33]&p[33]);
carry_out[34] = (g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))));
g[34] = a[34]&b_not[34];
p[34] = a[34]^b_not[34];

sum[34]= (p[34]^carry_in[34]);
carry_in[35] = (g[34]|carry_in[34]&p[34]);
carry_out[35] = (g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))));
g[35] = a[35]&b_not[35];
p[35] = a[35]^b_not[35];

sum[35]= (p[35]^carry_in[35]);
carry_in[36] = (g[35]|carry_in[35]&p[35]);
carry_out[36] = (g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))));
g[36] = a[36]&b_not[36];
p[36] = a[36]^b_not[36];

sum[36]= (p[36]^carry_in[36]);
carry_in[37] = (g[36]|carry_in[36]&p[36]);
carry_out[37] = (g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))));
g[37] = a[37]&b_not[37];
p[37] = a[37]^b_not[37];

sum[37]= (p[37]^carry_in[37]);
carry_in[38] = (g[37]|carry_in[37]&p[37]);
carry_out[38] = (g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))));
g[38] = a[38]&b_not[38];
p[38] = a[38]^b_not[38];

sum[38]= (p[38]^carry_in[38]);
carry_in[39] = (g[38]|carry_in[38]&p[38]);
carry_out[39] = (g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))));
g[39] = a[39]&b_not[39];
p[39] = a[39]^b_not[39];

sum[39]= (p[39]^carry_in[39]);
carry_in[40] = (g[39]|carry_in[39]&p[39]);
carry_out[40] = (g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))));
g[40] = a[40]&b_not[40];
p[40] = a[40]^b_not[40];

sum[40]= (p[40]^carry_in[40]);
carry_in[41] = (g[40]|carry_in[40]&p[40]);
carry_out[41] = (g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))));
g[41] = a[41]&b_not[41];
p[41] = a[41]^b_not[41];

sum[41]= (p[41]^carry_in[41]);
carry_in[42] = (g[41]|carry_in[41]&p[41]);
carry_out[42] = (g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))));
g[42] = a[42]&b_not[42];
p[42] = a[42]^b_not[42];

sum[42]= (p[42]^carry_in[42]);
carry_in[43] = (g[42]|carry_in[42]&p[42]);
carry_out[43] = (g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))));
g[43] = a[43]&b_not[43];
p[43] = a[43]^b_not[43];

sum[43]= (p[43]^carry_in[43]);
carry_in[44] = (g[43]|carry_in[43]&p[43]);
carry_out[44] = (g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))));
g[44] = a[44]&b_not[44];
p[44] = a[44]^b_not[44];

sum[44]= (p[44]^carry_in[44]);
carry_in[45] = (g[44]|carry_in[44]&p[44]);
carry_out[45] = (g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))));
g[45] = a[45]&b_not[45];
p[45] = a[45]^b_not[45];

sum[45]= (p[45]^carry_in[45]);
carry_in[46] = (g[45]|carry_in[45]&p[45]);
carry_out[46] = (g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))));
g[46] = a[46]&b_not[46];
p[46] = a[46]^b_not[46];

sum[46]= (p[46]^carry_in[46]);
carry_in[47] = (g[46]|carry_in[46]&p[46]);
carry_out[47] = (g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))));
g[47] = a[47]&b_not[47];
p[47] = a[47]^b_not[47];

sum[47]= (p[47]^carry_in[47]);
carry_in[48] = (g[47]|carry_in[47]&p[47]);
carry_out[48] = (g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))));
g[48] = a[48]&b_not[48];
p[48] = a[48]^b_not[48];

sum[48]= (p[48]^carry_in[48]);
carry_in[49] = (g[48]|carry_in[48]&p[48]);
carry_out[49] = (g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))));
g[49] = a[49]&b_not[49];
p[49] = a[49]^b_not[49];

sum[49]= (p[49]^carry_in[49]);
carry_in[50] = (g[49]|carry_in[49]&p[49]);
carry_out[50] = (g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))));
g[50] = a[50]&b_not[50];
p[50] = a[50]^b_not[50];

sum[50]= (p[50]^carry_in[50]);
carry_in[51] = (g[50]|carry_in[50]&p[50]);
carry_out[51] = (g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))));
g[51] = a[51]&b_not[51];
p[51] = a[51]^b_not[51];

sum[51]= (p[51]^carry_in[51]);
carry_in[52] = (g[51]|carry_in[51]&p[51]);
carry_out[52] = (g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))));
g[52] = a[52]&b_not[52];
p[52] = a[52]^b_not[52];

sum[52]= (p[52]^carry_in[52]);
carry_in[53] = (g[52]|carry_in[52]&p[52]);
carry_out[53] = (g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))));
g[53] = a[53]&b_not[53];
p[53] = a[53]^b_not[53];

sum[53]= (p[53]^carry_in[53]);
carry_in[54] = (g[53]|carry_in[53]&p[53]);
carry_out[54] = (g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[54] = a[54]&b_not[54];
p[54] = a[54]^b_not[54];

sum[54]= (p[54]^carry_in[54]);
carry_in[55] = (g[54]|carry_in[54]&p[54]);
carry_out[55] = (g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[55] = a[55]&b_not[55];
p[55] = a[55]^b_not[55];

sum[55]= (p[55]^carry_in[55]);
carry_in[56] = (g[55]|carry_in[55]&p[55]);
carry_out[56] = (g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[56] = a[56]&b_not[56];
p[56] = a[56]^b_not[56];

sum[56]= (p[56]^carry_in[56]);
carry_in[57] = (g[56]|carry_in[56]&p[56]);
carry_out[57] = (g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[57] = a[57]&b_not[57];
p[57] = a[57]^b_not[57];

sum[57]= (p[57]^carry_in[57]);
carry_in[58] = (g[57]|carry_in[57]&p[57]);
carry_out[58] = (g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[58] = a[58]&b_not[58];
p[58] = a[58]^b_not[58];

sum[58]= (p[58]^carry_in[58]);
carry_in[59] = (g[58]|carry_in[58]&p[58]);
carry_out[59] = (g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[59] = a[59]&b_not[59];
p[59] = a[59]^b_not[59];

sum[59]= (p[59]^carry_in[59]);
carry_in[60] = (g[59]|carry_in[59]&p[59]);
carry_out[60] = (g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[60] = a[60]&b_not[60];
p[60] = a[60]^b_not[60];

sum[60]= (p[60]^carry_in[60]);
carry_in[61] = (g[60]|carry_in[60]&p[60]);
carry_out[61] = (g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[61] = a[61]&b_not[61];
p[61] = a[61]^b_not[61];

sum[61]= (p[61]^carry_in[61]);
carry_in[62] = (g[61]|carry_in[61]&p[61]);
carry_out[62] = (g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[62] = a[62]&b_not[62];
p[62] = a[62]^b_not[62];

sum[62]= (p[62]^carry_in[62]);
carry_in[63] = (g[62]|carry_in[62]&p[62]);
carry_out[63] = (g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[63] = a[63]&b_not[63];
p[63] = a[63]^b_not[63];

sum[63]= (p[63]^carry_in[63]);
carry_in[64] = (g[63]|carry_in[63]&p[63]);
carry_out[64] = (g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[64] = a[64]&b_not[64];
p[64] = a[64]^b_not[64];

sum[64]= (p[64]^carry_in[64]);
carry_in[65] = (g[64]|carry_in[64]&p[64]);
carry_out[65] = (g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[65] = a[65]&b_not[65];
p[65] = a[65]^b_not[65];

sum[65]= (p[65]^carry_in[65]);
carry_in[66] = (g[65]|carry_in[65]&p[65]);
carry_out[66] = (g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[66] = a[66]&b_not[66];
p[66] = a[66]^b_not[66];

sum[66]= (p[66]^carry_in[66]);
carry_in[67] = (g[66]|carry_in[66]&p[66]);
carry_out[67] = (g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[67] = a[67]&b_not[67];
p[67] = a[67]^b_not[67];

sum[67]= (p[67]^carry_in[67]);
carry_in[68] = (g[67]|carry_in[67]&p[67]);
carry_out[68] = (g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[68] = a[68]&b_not[68];
p[68] = a[68]^b_not[68];

sum[68]= (p[68]^carry_in[68]);
carry_in[69] = (g[68]|carry_in[68]&p[68]);
carry_out[69] = (g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[69] = a[69]&b_not[69];
p[69] = a[69]^b_not[69];

sum[69]= (p[69]^carry_in[69]);
carry_in[70] = (g[69]|carry_in[69]&p[69]);
carry_out[70] = (g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[70] = a[70]&b_not[70];
p[70] = a[70]^b_not[70];

sum[70]= (p[70]^carry_in[70]);
carry_in[71] = (g[70]|carry_in[70]&p[70]);
carry_out[71] = (g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[71] = a[71]&b_not[71];
p[71] = a[71]^b_not[71];

sum[71]= (p[71]^carry_in[71]);
carry_in[72] = (g[71]|carry_in[71]&p[71]);
carry_out[72] = (g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[72] = a[72]&b_not[72];
p[72] = a[72]^b_not[72];

sum[72]= (p[72]^carry_in[72]);
carry_in[73] = (g[72]|carry_in[72]&p[72]);
carry_out[73] = (g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[73] = a[73]&b_not[73];
p[73] = a[73]^b_not[73];

sum[73]= (p[73]^carry_in[73]);
carry_in[74] = (g[73]|carry_in[73]&p[73]);
carry_out[74] = (g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[74] = a[74]&b_not[74];
p[74] = a[74]^b_not[74];

sum[74]= (p[74]^carry_in[74]);
carry_in[75] = (g[74]|carry_in[74]&p[74]);
carry_out[75] = (g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[75] = a[75]&b_not[75];
p[75] = a[75]^b_not[75];

sum[75]= (p[75]^carry_in[75]);
carry_in[76] = (g[75]|carry_in[75]&p[75]);
carry_out[76] = (g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[76] = a[76]&b_not[76];
p[76] = a[76]^b_not[76];

sum[76]= (p[76]^carry_in[76]);
carry_in[77] = (g[76]|carry_in[76]&p[76]);
carry_out[77] = (g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[77] = a[77]&b_not[77];
p[77] = a[77]^b_not[77];

sum[77]= (p[77]^carry_in[77]);
carry_in[78] = (g[77]|carry_in[77]&p[77]);
carry_out[78] = (g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[78] = a[78]&b_not[78];
p[78] = a[78]^b_not[78];

sum[78]= (p[78]^carry_in[78]);
carry_in[79] = (g[78]|carry_in[78]&p[78]);
carry_out[79] = (g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[79] = a[79]&b_not[79];
p[79] = a[79]^b_not[79];

sum[79]= (p[79]^carry_in[79]);
carry_in[80] = (g[79]|carry_in[79]&p[79]);
carry_out[80] = (g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[80] = a[80]&b_not[80];
p[80] = a[80]^b_not[80];

sum[80]= (p[80]^carry_in[80]);
carry_in[81] = (g[80]|carry_in[80]&p[80]);
carry_out[81] = (g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[81] = a[81]&b_not[81];
p[81] = a[81]^b_not[81];

sum[81]= (p[81]^carry_in[81]);
carry_in[82] = (g[81]|carry_in[81]&p[81]);
carry_out[82] = (g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[82] = a[82]&b_not[82];
p[82] = a[82]^b_not[82];

sum[82]= (p[82]^carry_in[82]);
carry_in[83] = (g[82]|carry_in[82]&p[82]);
carry_out[83] = (g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[83] = a[83]&b_not[83];
p[83] = a[83]^b_not[83];

sum[83]= (p[83]^carry_in[83]);
carry_in[84] = (g[83]|carry_in[83]&p[83]);
carry_out[84] = (g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[84] = a[84]&b_not[84];
p[84] = a[84]^b_not[84];

sum[84]= (p[84]^carry_in[84]);
carry_in[85] = (g[84]|carry_in[84]&p[84]);
carry_out[85] = (g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[85] = a[85]&b_not[85];
p[85] = a[85]^b_not[85];

sum[85]= (p[85]^carry_in[85]);
carry_in[86] = (g[85]|carry_in[85]&p[85]);
carry_out[86] = (g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[86] = a[86]&b_not[86];
p[86] = a[86]^b_not[86];

sum[86]= (p[86]^carry_in[86]);
carry_in[87] = (g[86]|carry_in[86]&p[86]);
carry_out[87] = (g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[87] = a[87]&b_not[87];
p[87] = a[87]^b_not[87];

sum[87]= (p[87]^carry_in[87]);
carry_in[88] = (g[87]|carry_in[87]&p[87]);
carry_out[88] = (g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[88] = a[88]&b_not[88];
p[88] = a[88]^b_not[88];

sum[88]= (p[88]^carry_in[88]);
carry_in[89] = (g[88]|carry_in[88]&p[88]);
carry_out[89] = (g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[89] = a[89]&b_not[89];
p[89] = a[89]^b_not[89];

sum[89]= (p[89]^carry_in[89]);
carry_in[90] = (g[89]|carry_in[89]&p[89]);
carry_out[90] = (g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[90] = a[90]&b_not[90];
p[90] = a[90]^b_not[90];

sum[90]= (p[90]^carry_in[90]);
carry_in[91] = (g[90]|carry_in[90]&p[90]);
carry_out[91] = (g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[91] = a[91]&b_not[91];
p[91] = a[91]^b_not[91];

sum[91]= (p[91]^carry_in[91]);
carry_in[92] = (g[91]|carry_in[91]&p[91]);
carry_out[92] = (g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[92] = a[92]&b_not[92];
p[92] = a[92]^b_not[92];

sum[92]= (p[92]^carry_in[92]);
carry_in[93] = (g[92]|carry_in[92]&p[92]);
carry_out[93] = (g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[93] = a[93]&b_not[93];
p[93] = a[93]^b_not[93];

sum[93]= (p[93]^carry_in[93]);
carry_in[94] = (g[93]|carry_in[93]&p[93]);
carry_out[94] = (g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[94] = a[94]&b_not[94];
p[94] = a[94]^b_not[94];

sum[94]= (p[94]^carry_in[94]);
carry_in[95] = (g[94]|carry_in[94]&p[94]);
carry_out[95] = (g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[95] = a[95]&b_not[95];
p[95] = a[95]^b_not[95];

sum[95]= (p[95]^carry_in[95]);
carry_in[96] = (g[95]|carry_in[95]&p[95]);
carry_out[96] = (g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[96] = a[96]&b_not[96];
p[96] = a[96]^b_not[96];

sum[96]= (p[96]^carry_in[96]);
carry_in[97] = (g[96]|carry_in[96]&p[96]);
carry_out[97] = (g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[97] = a[97]&b_not[97];
p[97] = a[97]^b_not[97];

sum[97]= (p[97]^carry_in[97]);
carry_in[98] = (g[97]|carry_in[97]&p[97]);
carry_out[98] = (g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[98] = a[98]&b_not[98];
p[98] = a[98]^b_not[98];

sum[98]= (p[98]^carry_in[98]);
carry_in[99] = (g[98]|carry_in[98]&p[98]);
carry_out[99] = (g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[99] = a[99]&b_not[99];
p[99] = a[99]^b_not[99];

sum[99]= (p[99]^carry_in[99]);
carry_in[100] = (g[99]|carry_in[99]&p[99]);
carry_out[100] = (g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[100] = a[100]&b_not[100];
p[100] = a[100]^b_not[100];

sum[100]= (p[100]^carry_in[100]);
carry_in[101] = (g[100]|carry_in[100]&p[100]);
carry_out[101] = (g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[101] = a[101]&b_not[101];
p[101] = a[101]^b_not[101];

sum[101]= (p[101]^carry_in[101]);
carry_in[102] = (g[101]|carry_in[101]&p[101]);
carry_out[102] = (g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[102] = a[102]&b_not[102];
p[102] = a[102]^b_not[102];

sum[102]= (p[102]^carry_in[102]);
carry_in[103] = (g[102]|carry_in[102]&p[102]);
carry_out[103] = (g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[103] = a[103]&b_not[103];
p[103] = a[103]^b_not[103];

sum[103]= (p[103]^carry_in[103]);
carry_in[104] = (g[103]|carry_in[103]&p[103]);
carry_out[104] = (g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[104] = a[104]&b_not[104];
p[104] = a[104]^b_not[104];

sum[104]= (p[104]^carry_in[104]);
carry_in[105] = (g[104]|carry_in[104]&p[104]);
carry_out[105] = (g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[105] = a[105]&b_not[105];
p[105] = a[105]^b_not[105];

sum[105]= (p[105]^carry_in[105]);
carry_in[106] = (g[105]|carry_in[105]&p[105]);
carry_out[106] = (g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[106] = a[106]&b_not[106];
p[106] = a[106]^b_not[106];

sum[106]= (p[106]^carry_in[106]);
carry_in[107] = (g[106]|carry_in[106]&p[106]);
carry_out[107] = (g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[107] = a[107]&b_not[107];
p[107] = a[107]^b_not[107];

sum[107]= (p[107]^carry_in[107]);
carry_in[108] = (g[107]|carry_in[107]&p[107]);
carry_out[108] = (g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[108] = a[108]&b_not[108];
p[108] = a[108]^b_not[108];

sum[108]= (p[108]^carry_in[108]);
carry_in[109] = (g[108]|carry_in[108]&p[108]);
carry_out[109] = (g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[109] = a[109]&b_not[109];
p[109] = a[109]^b_not[109];

sum[109]= (p[109]^carry_in[109]);
carry_in[110] = (g[109]|carry_in[109]&p[109]);
carry_out[110] = (g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[110] = a[110]&b_not[110];
p[110] = a[110]^b_not[110];

sum[110]= (p[110]^carry_in[110]);
carry_in[111] = (g[110]|carry_in[110]&p[110]);
carry_out[111] = (g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[111] = a[111]&b_not[111];
p[111] = a[111]^b_not[111];

sum[111]= (p[111]^carry_in[111]);
carry_in[112] = (g[111]|carry_in[111]&p[111]);
carry_out[112] = (g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[112] = a[112]&b_not[112];
p[112] = a[112]^b_not[112];

sum[112]= (p[112]^carry_in[112]);
carry_in[113] = (g[112]|carry_in[112]&p[112]);
carry_out[113] = (g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[113] = a[113]&b_not[113];
p[113] = a[113]^b_not[113];

sum[113]= (p[113]^carry_in[113]);
carry_in[114] = (g[113]|carry_in[113]&p[113]);
carry_out[114] = (g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[114] = a[114]&b_not[114];
p[114] = a[114]^b_not[114];

sum[114]= (p[114]^carry_in[114]);
carry_in[115] = (g[114]|carry_in[114]&p[114]);
carry_out[115] = (g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[115] = a[115]&b_not[115];
p[115] = a[115]^b_not[115];

sum[115]= (p[115]^carry_in[115]);
carry_in[116] = (g[115]|carry_in[115]&p[115]);
carry_out[116] = (g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[116] = a[116]&b_not[116];
p[116] = a[116]^b_not[116];

sum[116]= (p[116]^carry_in[116]);
carry_in[117] = (g[116]|carry_in[116]&p[116]);
carry_out[117] = (g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[117] = a[117]&b_not[117];
p[117] = a[117]^b_not[117];

sum[117]= (p[117]^carry_in[117]);
carry_in[118] = (g[117]|carry_in[117]&p[117]);
carry_out[118] = (g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[118] = a[118]&b_not[118];
p[118] = a[118]^b_not[118];

sum[118]= (p[118]^carry_in[118]);
carry_in[119] = (g[118]|carry_in[118]&p[118]);
carry_out[119] = (g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[119] = a[119]&b_not[119];
p[119] = a[119]^b_not[119];

sum[119]= (p[119]^carry_in[119]);
carry_in[120] = (g[119]|carry_in[119]&p[119]);
carry_out[120] = (g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[120] = a[120]&b_not[120];
p[120] = a[120]^b_not[120];

sum[120]= (p[120]^carry_in[120]);
carry_in[121] = (g[120]|carry_in[120]&p[120]);
carry_out[121] = (g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[121] = a[121]&b_not[121];
p[121] = a[121]^b_not[121];

sum[121]= (p[121]^carry_in[121]);
carry_in[122] = (g[121]|carry_in[121]&p[121]);
carry_out[122] = (g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[122] = a[122]&b_not[122];
p[122] = a[122]^b_not[122];

sum[122]= (p[122]^carry_in[122]);
carry_in[123] = (g[122]|carry_in[122]&p[122]);
carry_out[123] = (g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[123] = a[123]&b_not[123];
p[123] = a[123]^b_not[123];

sum[123]= (p[123]^carry_in[123]);
carry_in[124] = (g[123]|carry_in[123]&p[123]);
carry_out[124] = (g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[124] = a[124]&b_not[124];
p[124] = a[124]^b_not[124];

sum[124]= (p[124]^carry_in[124]);
carry_in[125] = (g[124]|carry_in[124]&p[124]);
carry_out[125] = (g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[125] = a[125]&b_not[125];
p[125] = a[125]^b_not[125];

sum[125]= (p[125]^carry_in[125]);
carry_in[126] = (g[125]|carry_in[125]&p[125]);
carry_out[126] = (g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[126] = a[126]&b_not[126];
p[126] = a[126]^b_not[126];

sum[126]= (p[126]^carry_in[126]);
carry_in[127] = (g[126]|carry_in[126]&p[126]);
carry_out[127] = (g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[127] = a[127]&b_not[127];
p[127] = a[127]^b_not[127];

sum[127]= (p[127]^carry_in[127]);
carry_in[128] = (g[127]|carry_in[127]&p[127]);
carry_out[128] = (g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[128] = a[128]&b_not[128];
p[128] = a[128]^b_not[128];

sum[128]= (p[128]^carry_in[128]);
carry_in[129] = (g[128]|carry_in[128]&p[128]);
carry_out[129] = (g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[129] = a[129]&b_not[129];
p[129] = a[129]^b_not[129];

sum[129]= (p[129]^carry_in[129]);
carry_in[130] = (g[129]|carry_in[129]&p[129]);
carry_out[130] = (g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[130] = a[130]&b_not[130];
p[130] = a[130]^b_not[130];

sum[130]= (p[130]^carry_in[130]);
carry_in[131] = (g[130]|carry_in[130]&p[130]);
carry_out[131] = (g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[131] = a[131]&b_not[131];
p[131] = a[131]^b_not[131];

sum[131]= (p[131]^carry_in[131]);
carry_in[132] = (g[131]|carry_in[131]&p[131]);
carry_out[132] = (g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[132] = a[132]&b_not[132];
p[132] = a[132]^b_not[132];

sum[132]= (p[132]^carry_in[132]);
carry_in[133] = (g[132]|carry_in[132]&p[132]);
carry_out[133] = (g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[133] = a[133]&b_not[133];
p[133] = a[133]^b_not[133];

sum[133]= (p[133]^carry_in[133]);
carry_in[134] = (g[133]|carry_in[133]&p[133]);
carry_out[134] = (g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[134] = a[134]&b_not[134];
p[134] = a[134]^b_not[134];

sum[134]= (p[134]^carry_in[134]);
carry_in[135] = (g[134]|carry_in[134]&p[134]);
carry_out[135] = (g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[135] = a[135]&b_not[135];
p[135] = a[135]^b_not[135];

sum[135]= (p[135]^carry_in[135]);
carry_in[136] = (g[135]|carry_in[135]&p[135]);
carry_out[136] = (g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[136] = a[136]&b_not[136];
p[136] = a[136]^b_not[136];

sum[136]= (p[136]^carry_in[136]);
carry_in[137] = (g[136]|carry_in[136]&p[136]);
carry_out[137] = (g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[137] = a[137]&b_not[137];
p[137] = a[137]^b_not[137];

sum[137]= (p[137]^carry_in[137]);
carry_in[138] = (g[137]|carry_in[137]&p[137]);
carry_out[138] = (g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[138] = a[138]&b_not[138];
p[138] = a[138]^b_not[138];

sum[138]= (p[138]^carry_in[138]);
carry_in[139] = (g[138]|carry_in[138]&p[138]);
carry_out[139] = (g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[139] = a[139]&b_not[139];
p[139] = a[139]^b_not[139];

sum[139]= (p[139]^carry_in[139]);
carry_in[140] = (g[139]|carry_in[139]&p[139]);
carry_out[140] = (g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[140] = a[140]&b_not[140];
p[140] = a[140]^b_not[140];

sum[140]= (p[140]^carry_in[140]);
carry_in[141] = (g[140]|carry_in[140]&p[140]);
carry_out[141] = (g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[141] = a[141]&b_not[141];
p[141] = a[141]^b_not[141];

sum[141]= (p[141]^carry_in[141]);
carry_in[142] = (g[141]|carry_in[141]&p[141]);
carry_out[142] = (g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[142] = a[142]&b_not[142];
p[142] = a[142]^b_not[142];

sum[142]= (p[142]^carry_in[142]);
carry_in[143] = (g[142]|carry_in[142]&p[142]);
carry_out[143] = (g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[143] = a[143]&b_not[143];
p[143] = a[143]^b_not[143];

sum[143]= (p[143]^carry_in[143]);
carry_in[144] = (g[143]|carry_in[143]&p[143]);
carry_out[144] = (g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[144] = a[144]&b_not[144];
p[144] = a[144]^b_not[144];

sum[144]= (p[144]^carry_in[144]);
carry_in[145] = (g[144]|carry_in[144]&p[144]);
carry_out[145] = (g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[145] = a[145]&b_not[145];
p[145] = a[145]^b_not[145];

sum[145]= (p[145]^carry_in[145]);
carry_in[146] = (g[145]|carry_in[145]&p[145]);
carry_out[146] = (g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[146] = a[146]&b_not[146];
p[146] = a[146]^b_not[146];

sum[146]= (p[146]^carry_in[146]);
carry_in[147] = (g[146]|carry_in[146]&p[146]);
carry_out[147] = (g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[147] = a[147]&b_not[147];
p[147] = a[147]^b_not[147];

sum[147]= (p[147]^carry_in[147]);
carry_in[148] = (g[147]|carry_in[147]&p[147]);
carry_out[148] = (g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[148] = a[148]&b_not[148];
p[148] = a[148]^b_not[148];

sum[148]= (p[148]^carry_in[148]);
carry_in[149] = (g[148]|carry_in[148]&p[148]);
carry_out[149] = (g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[149] = a[149]&b_not[149];
p[149] = a[149]^b_not[149];

sum[149]= (p[149]^carry_in[149]);
carry_in[150] = (g[149]|carry_in[149]&p[149]);
carry_out[150] = (g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[150] = a[150]&b_not[150];
p[150] = a[150]^b_not[150];

sum[150]= (p[150]^carry_in[150]);
carry_in[151] = (g[150]|carry_in[150]&p[150]);
carry_out[151] = (g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[151] = a[151]&b_not[151];
p[151] = a[151]^b_not[151];

sum[151]= (p[151]^carry_in[151]);
carry_in[152] = (g[151]|carry_in[151]&p[151]);
carry_out[152] = (g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[152] = a[152]&b_not[152];
p[152] = a[152]^b_not[152];

sum[152]= (p[152]^carry_in[152]);
carry_in[153] = (g[152]|carry_in[152]&p[152]);
carry_out[153] = (g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[153] = a[153]&b_not[153];
p[153] = a[153]^b_not[153];

sum[153]= (p[153]^carry_in[153]);
carry_in[154] = (g[153]|carry_in[153]&p[153]);
carry_out[154] = (g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[154] = a[154]&b_not[154];
p[154] = a[154]^b_not[154];

sum[154]= (p[154]^carry_in[154]);
carry_in[155] = (g[154]|carry_in[154]&p[154]);
carry_out[155] = (g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[155] = a[155]&b_not[155];
p[155] = a[155]^b_not[155];

sum[155]= (p[155]^carry_in[155]);
carry_in[156] = (g[155]|carry_in[155]&p[155]);
carry_out[156] = (g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[156] = a[156]&b_not[156];
p[156] = a[156]^b_not[156];

sum[156]= (p[156]^carry_in[156]);
carry_in[157] = (g[156]|carry_in[156]&p[156]);
carry_out[157] = (g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[157] = a[157]&b_not[157];
p[157] = a[157]^b_not[157];

sum[157]= (p[157]^carry_in[157]);
carry_in[158] = (g[157]|carry_in[157]&p[157]);
carry_out[158] = (g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[158] = a[158]&b_not[158];
p[158] = a[158]^b_not[158];

sum[158]= (p[158]^carry_in[158]);
carry_in[159] = (g[158]|carry_in[158]&p[158]);
carry_out[159] = (g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[159] = a[159]&b_not[159];
p[159] = a[159]^b_not[159];

sum[159]= (p[159]^carry_in[159]);
carry_in[160] = (g[159]|carry_in[159]&p[159]);
carry_out[160] = (g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[160] = a[160]&b_not[160];
p[160] = a[160]^b_not[160];

sum[160]= (p[160]^carry_in[160]);
carry_in[161] = (g[160]|carry_in[160]&p[160]);
carry_out[161] = (g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[161] = a[161]&b_not[161];
p[161] = a[161]^b_not[161];

sum[161]= (p[161]^carry_in[161]);
carry_in[162] = (g[161]|carry_in[161]&p[161]);
carry_out[162] = (g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[162] = a[162]&b_not[162];
p[162] = a[162]^b_not[162];

sum[162]= (p[162]^carry_in[162]);
carry_in[163] = (g[162]|carry_in[162]&p[162]);
carry_out[163] = (g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[163] = a[163]&b_not[163];
p[163] = a[163]^b_not[163];

sum[163]= (p[163]^carry_in[163]);
carry_in[164] = (g[163]|carry_in[163]&p[163]);
carry_out[164] = (g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[164] = a[164]&b_not[164];
p[164] = a[164]^b_not[164];

sum[164]= (p[164]^carry_in[164]);
carry_in[165] = (g[164]|carry_in[164]&p[164]);
carry_out[165] = (g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[165] = a[165]&b_not[165];
p[165] = a[165]^b_not[165];

sum[165]= (p[165]^carry_in[165]);
carry_in[166] = (g[165]|carry_in[165]&p[165]);
carry_out[166] = (g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[166] = a[166]&b_not[166];
p[166] = a[166]^b_not[166];

sum[166]= (p[166]^carry_in[166]);
carry_in[167] = (g[166]|carry_in[166]&p[166]);
carry_out[167] = (g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[167] = a[167]&b_not[167];
p[167] = a[167]^b_not[167];

sum[167]= (p[167]^carry_in[167]);
carry_in[168] = (g[167]|carry_in[167]&p[167]);
carry_out[168] = (g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[168] = a[168]&b_not[168];
p[168] = a[168]^b_not[168];

sum[168]= (p[168]^carry_in[168]);
carry_in[169] = (g[168]|carry_in[168]&p[168]);
carry_out[169] = (g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[169] = a[169]&b_not[169];
p[169] = a[169]^b_not[169];

sum[169]= (p[169]^carry_in[169]);
carry_in[170] = (g[169]|carry_in[169]&p[169]);
carry_out[170] = (g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[170] = a[170]&b_not[170];
p[170] = a[170]^b_not[170];

sum[170]= (p[170]^carry_in[170]);
carry_in[171] = (g[170]|carry_in[170]&p[170]);
carry_out[171] = (g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[171] = a[171]&b_not[171];
p[171] = a[171]^b_not[171];

sum[171]= (p[171]^carry_in[171]);
carry_in[172] = (g[171]|carry_in[171]&p[171]);
carry_out[172] = (g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[172] = a[172]&b_not[172];
p[172] = a[172]^b_not[172];

sum[172]= (p[172]^carry_in[172]);
carry_in[173] = (g[172]|carry_in[172]&p[172]);
carry_out[173] = (g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[173] = a[173]&b_not[173];
p[173] = a[173]^b_not[173];

sum[173]= (p[173]^carry_in[173]);
carry_in[174] = (g[173]|carry_in[173]&p[173]);
carry_out[174] = (g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[174] = a[174]&b_not[174];
p[174] = a[174]^b_not[174];

sum[174]= (p[174]^carry_in[174]);
carry_in[175] = (g[174]|carry_in[174]&p[174]);
carry_out[175] = (g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[175] = a[175]&b_not[175];
p[175] = a[175]^b_not[175];

sum[175]= (p[175]^carry_in[175]);
carry_in[176] = (g[175]|carry_in[175]&p[175]);
carry_out[176] = (g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[176] = a[176]&b_not[176];
p[176] = a[176]^b_not[176];

sum[176]= (p[176]^carry_in[176]);
carry_in[177] = (g[176]|carry_in[176]&p[176]);
carry_out[177] = (g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[177] = a[177]&b_not[177];
p[177] = a[177]^b_not[177];

sum[177]= (p[177]^carry_in[177]);
carry_in[178] = (g[177]|carry_in[177]&p[177]);
carry_out[178] = (g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[178] = a[178]&b_not[178];
p[178] = a[178]^b_not[178];

sum[178]= (p[178]^carry_in[178]);
carry_in[179] = (g[178]|carry_in[178]&p[178]);
carry_out[179] = (g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[179] = a[179]&b_not[179];
p[179] = a[179]^b_not[179];

sum[179]= (p[179]^carry_in[179]);
carry_in[180] = (g[179]|carry_in[179]&p[179]);
carry_out[180] = (g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[180] = a[180]&b_not[180];
p[180] = a[180]^b_not[180];

sum[180]= (p[180]^carry_in[180]);
carry_in[181] = (g[180]|carry_in[180]&p[180]);
carry_out[181] = (g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[181] = a[181]&b_not[181];
p[181] = a[181]^b_not[181];

sum[181]= (p[181]^carry_in[181]);
carry_in[182] = (g[181]|carry_in[181]&p[181]);
carry_out[182] = (g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[182] = a[182]&b_not[182];
p[182] = a[182]^b_not[182];

sum[182]= (p[182]^carry_in[182]);
carry_in[183] = (g[182]|carry_in[182]&p[182]);
carry_out[183] = (g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[183] = a[183]&b_not[183];
p[183] = a[183]^b_not[183];

sum[183]= (p[183]^carry_in[183]);
carry_in[184] = (g[183]|carry_in[183]&p[183]);
carry_out[184] = (g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[184] = a[184]&b_not[184];
p[184] = a[184]^b_not[184];

sum[184]= (p[184]^carry_in[184]);
carry_in[185] = (g[184]|carry_in[184]&p[184]);
carry_out[185] = (g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[185] = a[185]&b_not[185];
p[185] = a[185]^b_not[185];

sum[185]= (p[185]^carry_in[185]);
carry_in[186] = (g[185]|carry_in[185]&p[185]);
carry_out[186] = (g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[186] = a[186]&b_not[186];
p[186] = a[186]^b_not[186];

sum[186]= (p[186]^carry_in[186]);
carry_in[187] = (g[186]|carry_in[186]&p[186]);
carry_out[187] = (g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[187] = a[187]&b_not[187];
p[187] = a[187]^b_not[187];

sum[187]= (p[187]^carry_in[187]);
carry_in[188] = (g[187]|carry_in[187]&p[187]);
carry_out[188] = (g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[188] = a[188]&b_not[188];
p[188] = a[188]^b_not[188];

sum[188]= (p[188]^carry_in[188]);
carry_in[189] = (g[188]|carry_in[188]&p[188]);
carry_out[189] = (g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[189] = a[189]&b_not[189];
p[189] = a[189]^b_not[189];

sum[189]= (p[189]^carry_in[189]);
carry_in[190] = (g[189]|carry_in[189]&p[189]);
carry_out[190] = (g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[190] = a[190]&b_not[190];
p[190] = a[190]^b_not[190];

sum[190]= (p[190]^carry_in[190]);
carry_in[191] = (g[190]|carry_in[190]&p[190]);
carry_out[191] = (g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[191] = a[191]&b_not[191];
p[191] = a[191]^b_not[191];

sum[191]= (p[191]^carry_in[191]);
carry_in[192] = (g[191]|carry_in[191]&p[191]);
carry_out[192] = (g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[192] = a[192]&b_not[192];
p[192] = a[192]^b_not[192];

sum[192]= (p[192]^carry_in[192]);
carry_in[193] = (g[192]|carry_in[192]&p[192]);
carry_out[193] = (g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[193] = a[193]&b_not[193];
p[193] = a[193]^b_not[193];

sum[193]= (p[193]^carry_in[193]);
carry_in[194] = (g[193]|carry_in[193]&p[193]);
carry_out[194] = (g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[194] = a[194]&b_not[194];
p[194] = a[194]^b_not[194];

sum[194]= (p[194]^carry_in[194]);
carry_in[195] = (g[194]|carry_in[194]&p[194]);
carry_out[195] = (g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[195] = a[195]&b_not[195];
p[195] = a[195]^b_not[195];

sum[195]= (p[195]^carry_in[195]);
carry_in[196] = (g[195]|carry_in[195]&p[195]);
carry_out[196] = (g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[196] = a[196]&b_not[196];
p[196] = a[196]^b_not[196];

sum[196]= (p[196]^carry_in[196]);
carry_in[197] = (g[196]|carry_in[196]&p[196]);
carry_out[197] = (g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[197] = a[197]&b_not[197];
p[197] = a[197]^b_not[197];

sum[197]= (p[197]^carry_in[197]);
carry_in[198] = (g[197]|carry_in[197]&p[197]);
carry_out[198] = (g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[198] = a[198]&b_not[198];
p[198] = a[198]^b_not[198];

sum[198]= (p[198]^carry_in[198]);
carry_in[199] = (g[198]|carry_in[198]&p[198]);
carry_out[199] = (g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[199] = a[199]&b_not[199];
p[199] = a[199]^b_not[199];

sum[199]= (p[199]^carry_in[199]);
carry_in[200] = (g[199]|carry_in[199]&p[199]);
carry_out[200] = (g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[200] = a[200]&b_not[200];
p[200] = a[200]^b_not[200];

sum[200]= (p[200]^carry_in[200]);
carry_in[201] = (g[200]|carry_in[200]&p[200]);
carry_out[201] = (g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[201] = a[201]&b_not[201];
p[201] = a[201]^b_not[201];

sum[201]= (p[201]^carry_in[201]);
carry_in[202] = (g[201]|carry_in[201]&p[201]);
carry_out[202] = (g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[202] = a[202]&b_not[202];
p[202] = a[202]^b_not[202];

sum[202]= (p[202]^carry_in[202]);
carry_in[203] = (g[202]|carry_in[202]&p[202]);
carry_out[203] = (g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[203] = a[203]&b_not[203];
p[203] = a[203]^b_not[203];

sum[203]= (p[203]^carry_in[203]);
carry_in[204] = (g[203]|carry_in[203]&p[203]);
carry_out[204] = (g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[204] = a[204]&b_not[204];
p[204] = a[204]^b_not[204];

sum[204]= (p[204]^carry_in[204]);
carry_in[205] = (g[204]|carry_in[204]&p[204]);
carry_out[205] = (g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[205] = a[205]&b_not[205];
p[205] = a[205]^b_not[205];

sum[205]= (p[205]^carry_in[205]);
carry_in[206] = (g[205]|carry_in[205]&p[205]);
carry_out[206] = (g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[206] = a[206]&b_not[206];
p[206] = a[206]^b_not[206];

sum[206]= (p[206]^carry_in[206]);
carry_in[207] = (g[206]|carry_in[206]&p[206]);
carry_out[207] = (g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[207] = a[207]&b_not[207];
p[207] = a[207]^b_not[207];

sum[207]= (p[207]^carry_in[207]);
carry_in[208] = (g[207]|carry_in[207]&p[207]);
carry_out[208] = (g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[208] = a[208]&b_not[208];
p[208] = a[208]^b_not[208];

sum[208]= (p[208]^carry_in[208]);
carry_in[209] = (g[208]|carry_in[208]&p[208]);
carry_out[209] = (g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[209] = a[209]&b_not[209];
p[209] = a[209]^b_not[209];

sum[209]= (p[209]^carry_in[209]);
carry_in[210] = (g[209]|carry_in[209]&p[209]);
carry_out[210] = (g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[210] = a[210]&b_not[210];
p[210] = a[210]^b_not[210];

sum[210]= (p[210]^carry_in[210]);
carry_in[211] = (g[210]|carry_in[210]&p[210]);
carry_out[211] = (g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[211] = a[211]&b_not[211];
p[211] = a[211]^b_not[211];

sum[211]= (p[211]^carry_in[211]);
carry_in[212] = (g[211]|carry_in[211]&p[211]);
carry_out[212] = (g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[212] = a[212]&b_not[212];
p[212] = a[212]^b_not[212];

sum[212]= (p[212]^carry_in[212]);
carry_in[213] = (g[212]|carry_in[212]&p[212]);
carry_out[213] = (g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[213] = a[213]&b_not[213];
p[213] = a[213]^b_not[213];

sum[213]= (p[213]^carry_in[213]);
carry_in[214] = (g[213]|carry_in[213]&p[213]);
carry_out[214] = (g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[214] = a[214]&b_not[214];
p[214] = a[214]^b_not[214];

sum[214]= (p[214]^carry_in[214]);
carry_in[215] = (g[214]|carry_in[214]&p[214]);
carry_out[215] = (g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[215] = a[215]&b_not[215];
p[215] = a[215]^b_not[215];

sum[215]= (p[215]^carry_in[215]);
carry_in[216] = (g[215]|carry_in[215]&p[215]);
carry_out[216] = (g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[216] = a[216]&b_not[216];
p[216] = a[216]^b_not[216];

sum[216]= (p[216]^carry_in[216]);
carry_in[217] = (g[216]|carry_in[216]&p[216]);
carry_out[217] = (g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[217] = a[217]&b_not[217];
p[217] = a[217]^b_not[217];

sum[217]= (p[217]^carry_in[217]);
carry_in[218] = (g[217]|carry_in[217]&p[217]);
carry_out[218] = (g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[218] = a[218]&b_not[218];
p[218] = a[218]^b_not[218];

sum[218]= (p[218]^carry_in[218]);
carry_in[219] = (g[218]|carry_in[218]&p[218]);
carry_out[219] = (g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[219] = a[219]&b_not[219];
p[219] = a[219]^b_not[219];

sum[219]= (p[219]^carry_in[219]);
carry_in[220] = (g[219]|carry_in[219]&p[219]);
carry_out[220] = (g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[220] = a[220]&b_not[220];
p[220] = a[220]^b_not[220];

sum[220]= (p[220]^carry_in[220]);
carry_in[221] = (g[220]|carry_in[220]&p[220]);
carry_out[221] = (g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[221] = a[221]&b_not[221];
p[221] = a[221]^b_not[221];

sum[221]= (p[221]^carry_in[221]);
carry_in[222] = (g[221]|carry_in[221]&p[221]);
carry_out[222] = (g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[222] = a[222]&b_not[222];
p[222] = a[222]^b_not[222];

sum[222]= (p[222]^carry_in[222]);
carry_in[223] = (g[222]|carry_in[222]&p[222]);
carry_out[223] = (g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[223] = a[223]&b_not[223];
p[223] = a[223]^b_not[223];

sum[223]= (p[223]^carry_in[223]);
carry_in[224] = (g[223]|carry_in[223]&p[223]);
carry_out[224] = (g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[224] = a[224]&b_not[224];
p[224] = a[224]^b_not[224];

sum[224]= (p[224]^carry_in[224]);
carry_in[225] = (g[224]|carry_in[224]&p[224]);
carry_out[225] = (g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[225] = a[225]&b_not[225];
p[225] = a[225]^b_not[225];

sum[225]= (p[225]^carry_in[225]);
carry_in[226] = (g[225]|carry_in[225]&p[225]);
carry_out[226] = (g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[226] = a[226]&b_not[226];
p[226] = a[226]^b_not[226];

sum[226]= (p[226]^carry_in[226]);
carry_in[227] = (g[226]|carry_in[226]&p[226]);
carry_out[227] = (g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[227] = a[227]&b_not[227];
p[227] = a[227]^b_not[227];

sum[227]= (p[227]^carry_in[227]);
carry_in[228] = (g[227]|carry_in[227]&p[227]);
carry_out[228] = (g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[228] = a[228]&b_not[228];
p[228] = a[228]^b_not[228];

sum[228]= (p[228]^carry_in[228]);
carry_in[229] = (g[228]|carry_in[228]&p[228]);
carry_out[229] = (g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[229] = a[229]&b_not[229];
p[229] = a[229]^b_not[229];

sum[229]= (p[229]^carry_in[229]);
carry_in[230] = (g[229]|carry_in[229]&p[229]);
carry_out[230] = (g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[230] = a[230]&b_not[230];
p[230] = a[230]^b_not[230];

sum[230]= (p[230]^carry_in[230]);
carry_in[231] = (g[230]|carry_in[230]&p[230]);
carry_out[231] = (g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[231] = a[231]&b_not[231];
p[231] = a[231]^b_not[231];

sum[231]= (p[231]^carry_in[231]);
carry_in[232] = (g[231]|carry_in[231]&p[231]);
carry_out[232] = (g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[232] = a[232]&b_not[232];
p[232] = a[232]^b_not[232];

sum[232]= (p[232]^carry_in[232]);
carry_in[233] = (g[232]|carry_in[232]&p[232]);
carry_out[233] = (g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[233] = a[233]&b_not[233];
p[233] = a[233]^b_not[233];

sum[233]= (p[233]^carry_in[233]);
carry_in[234] = (g[233]|carry_in[233]&p[233]);
carry_out[234] = (g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[234] = a[234]&b_not[234];
p[234] = a[234]^b_not[234];

sum[234]= (p[234]^carry_in[234]);
carry_in[235] = (g[234]|carry_in[234]&p[234]);
carry_out[235] = (g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[235] = a[235]&b_not[235];
p[235] = a[235]^b_not[235];

sum[235]= (p[235]^carry_in[235]);
carry_in[236] = (g[235]|carry_in[235]&p[235]);
carry_out[236] = (g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[236] = a[236]&b_not[236];
p[236] = a[236]^b_not[236];

sum[236]= (p[236]^carry_in[236]);
carry_in[237] = (g[236]|carry_in[236]&p[236]);
carry_out[237] = (g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[237] = a[237]&b_not[237];
p[237] = a[237]^b_not[237];

sum[237]= (p[237]^carry_in[237]);
carry_in[238] = (g[237]|carry_in[237]&p[237]);
carry_out[238] = (g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[238] = a[238]&b_not[238];
p[238] = a[238]^b_not[238];

sum[238]= (p[238]^carry_in[238]);
carry_in[239] = (g[238]|carry_in[238]&p[238]);
carry_out[239] = (g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[239] = a[239]&b_not[239];
p[239] = a[239]^b_not[239];

sum[239]= (p[239]^carry_in[239]);
carry_in[240] = (g[239]|carry_in[239]&p[239]);
carry_out[240] = (g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[240] = a[240]&b_not[240];
p[240] = a[240]^b_not[240];

sum[240]= (p[240]^carry_in[240]);
carry_in[241] = (g[240]|carry_in[240]&p[240]);
carry_out[241] = (g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[241] = a[241]&b_not[241];
p[241] = a[241]^b_not[241];

sum[241]= (p[241]^carry_in[241]);
carry_in[242] = (g[241]|carry_in[241]&p[241]);
carry_out[242] = (g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[242] = a[242]&b_not[242];
p[242] = a[242]^b_not[242];

sum[242]= (p[242]^carry_in[242]);
carry_in[243] = (g[242]|carry_in[242]&p[242]);
carry_out[243] = (g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[243] = a[243]&b_not[243];
p[243] = a[243]^b_not[243];

sum[243]= (p[243]^carry_in[243]);
carry_in[244] = (g[243]|carry_in[243]&p[243]);
carry_out[244] = (g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[244] = a[244]&b_not[244];
p[244] = a[244]^b_not[244];

sum[244]= (p[244]^carry_in[244]);
carry_in[245] = (g[244]|carry_in[244]&p[244]);
carry_out[245] = (g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[245] = a[245]&b_not[245];
p[245] = a[245]^b_not[245];

sum[245]= (p[245]^carry_in[245]);
carry_in[246] = (g[245]|carry_in[245]&p[245]);
carry_out[246] = (g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[246] = a[246]&b_not[246];
p[246] = a[246]^b_not[246];

sum[246]= (p[246]^carry_in[246]);
carry_in[247] = (g[246]|carry_in[246]&p[246]);
carry_out[247] = (g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[247] = a[247]&b_not[247];
p[247] = a[247]^b_not[247];

sum[247]= (p[247]^carry_in[247]);
carry_in[248] = (g[247]|carry_in[247]&p[247]);
carry_out[248] = (g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[248] = a[248]&b_not[248];
p[248] = a[248]^b_not[248];

sum[248]= (p[248]^carry_in[248]);
carry_in[249] = (g[248]|carry_in[248]&p[248]);
carry_out[249] = (g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[249] = a[249]&b_not[249];
p[249] = a[249]^b_not[249];

sum[249]= (p[249]^carry_in[249]);
carry_in[250] = (g[249]|carry_in[249]&p[249]);
carry_out[250] = (g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[250] = a[250]&b_not[250];
p[250] = a[250]^b_not[250];

sum[250]= (p[250]^carry_in[250]);
carry_in[251] = (g[250]|carry_in[250]&p[250]);
carry_out[251] = (g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[251] = a[251]&b_not[251];
p[251] = a[251]^b_not[251];

sum[251]= (p[251]^carry_in[251]);
carry_in[252] = (g[251]|carry_in[251]&p[251]);
carry_out[252] = (g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[252] = a[252]&b_not[252];
p[252] = a[252]^b_not[252];

sum[252]= (p[252]^carry_in[252]);
carry_in[253] = (g[252]|carry_in[252]&p[252]);
carry_out[253] = (g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[253] = a[253]&b_not[253];
p[253] = a[253]^b_not[253];

sum[253]= (p[253]^carry_in[253]);
carry_in[254] = (g[253]|carry_in[253]&p[253]);
carry_out[254] = (g[253] | p[253] &(g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[254] = a[254]&b_not[254];
p[254] = a[254]^b_not[254];

sum[254]= (p[254]^carry_in[254]);
carry_in[255] = (g[254]|carry_in[254]&p[254]);
carry_out[255] = (g[254] | p[254] &(g[253] | p[253] &(g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


g[255] = a[255]&b_not[255];
p[255] = a[255]^b_not[255];
sum[255] = (p[255]^carry_in[255]);
carry_out_overflow = (g[255] | p[255] & (g[254] | p[254] &(g[253] | p[253] &(g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


end
endmodule
