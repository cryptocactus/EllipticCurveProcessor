module P_Rom (
				output signed [255:0]P_Rom_const,
				output signed [255:0]B_Rom_const,
				output signed [255:0]A_Rom_const,
				output carry_in_n,
				output carry_in_2
);

assign A_Rom_const = 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798;
assign P_Rom_const = 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f;
assign B_Rom_const = 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8;
assign carry_in_n = 1'b0;
assign carry_in_2 = 1'b1;

endmodule
