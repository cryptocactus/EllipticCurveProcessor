//256-bit Carry Look Ahead Adder with overflow bit
//Created by: Colter Sisler, Scott Everitt, Steven Dougherty
//Team: Nighthawk
//Rev: 3.0
//2-22-2017


module adder_256 (
  input signed [255:0] a,
  input signed [255:0] b,
  input carry_in_n,
  output reg signed [255:0] sum,
  output reg carry_out_overflow
);


reg signed [255:0] g,p;
reg signed [255:0] carry_in;
reg signed [255:0] carry_out;

always @* begin


 #0


carry_out[1] = (((a[0]^b[0])&carry_in_n)|(a[0]&b[0]));
g[0] = a[0]&b[0];
p[0] = a[0]^b[0];
sum[0] = p[0]^carry_in_n;
carry_in[0] = carry_in_n;
carry_in[1] = (g[0] | carry_in[0]&p[0]);

g[1] = a[1]&b[1];
p[1] = a[1]^b[1];
sum[1]= (p[1]^carry_in[1]);
carry_in[2] = (g[1]|carry_in[1]&p[1]);
carry_out[2] = (g[1] | p[1] &(g[0] | carry_in[0]&p[0]));

g[2] = a[2]&b[2];
p[2] = a[2]^b[2];
sum[2]= (p[2]^carry_in[2]);
carry_in[3] = (g[2]|carry_in[2]&p[2]);
carry_out[3] = (g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])));

g[3] = a[3]&b[3];
p[3] = a[3]^b[3];
sum[3]= (p[3]^carry_in[3]);
carry_in[4] = (g[3]|carry_in[3]&p[3]);
carry_out[4] = (g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))));
g[4] = a[4]&b[4];
p[4] = a[4]^b[4];

sum[4]= (p[4]^carry_in[4]);
carry_in[5] = (g[4]|carry_in[4]&p[4]);
carry_out[5] = (g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))));
g[5] = a[5]&b[5];
p[5] = a[5]^b[5];

sum[5]= (p[5]^carry_in[5]);
carry_in[6] = (g[5]|carry_in[5]&p[5]);
carry_out[6] = (g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))));
g[6] = a[6]&b[6];
p[6] = a[6]^b[6];

sum[6]= (p[6]^carry_in[6]);
carry_in[7] = (g[6]|carry_in[6]&p[6]);
carry_out[7] = (g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))));
g[7] = a[7]&b[7];
p[7] = a[7]^b[7];

sum[7]= (p[7]^carry_in[7]);
carry_in[8] = (g[7]|carry_in[7]&p[7]);
carry_out[8] = (g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))));
g[8] = a[8]&b[8];
p[8] = a[8]^b[8];

sum[8]= (p[8]^carry_in[8]);
carry_in[9] = (g[8]|carry_in[8]&p[8]);
carry_out[9] = (g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))));
g[9] = a[9]&b[9];
p[9] = a[9]^b[9];

sum[9]= (p[9]^carry_in[9]);
carry_in[10] = (g[9]|carry_in[9]&p[9]);
carry_out[10] = (g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))));
g[10] = a[10]&b[10];
p[10] = a[10]^b[10];

sum[10]= (p[10]^carry_in[10]);
carry_in[11] = (g[10]|carry_in[10]&p[10]);
carry_out[11] = (g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))));
g[11] = a[11]&b[11];
p[11] = a[11]^b[11];

sum[11]= (p[11]^carry_in[11]);
carry_in[12] = (g[11]|carry_in[11]&p[11]);
carry_out[12] = (g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))));
g[12] = a[12]&b[12];
p[12] = a[12]^b[12];

sum[12]= (p[12]^carry_in[12]);
carry_in[13] = (g[12]|carry_in[12]&p[12]);
carry_out[13] = (g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))));
g[13] = a[13]&b[13];
p[13] = a[13]^b[13];

sum[13]= (p[13]^carry_in[13]);
carry_in[14] = (g[13]|carry_in[13]&p[13]);
carry_out[14] = (g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))));
g[14] = a[14]&b[14];
p[14] = a[14]^b[14];

sum[14]= (p[14]^carry_in[14]);
carry_in[15] = (g[14]|carry_in[14]&p[14]);
carry_out[15] = (g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))));
g[15] = a[15]&b[15];
p[15] = a[15]^b[15];

sum[15]= (p[15]^carry_in[15]);
carry_in[16] = (g[15]|carry_in[15]&p[15]);
carry_out[16] = (g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))));
g[16] = a[16]&b[16];
p[16] = a[16]^b[16];

sum[16]= (p[16]^carry_in[16]);
carry_in[17] = (g[16]|carry_in[16]&p[16]);
carry_out[17] = (g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))));
g[17] = a[17]&b[17];
p[17] = a[17]^b[17];

sum[17]= (p[17]^carry_in[17]);
carry_in[18] = (g[17]|carry_in[17]&p[17]);
carry_out[18] = (g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))));
g[18] = a[18]&b[18];
p[18] = a[18]^b[18];

sum[18]= (p[18]^carry_in[18]);
carry_in[19] = (g[18]|carry_in[18]&p[18]);
carry_out[19] = (g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))));
g[19] = a[19]&b[19];
p[19] = a[19]^b[19];

sum[19]= (p[19]^carry_in[19]);
carry_in[20] = (g[19]|carry_in[19]&p[19]);
carry_out[20] = (g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))));
g[20] = a[20]&b[20];
p[20] = a[20]^b[20];

sum[20]= (p[20]^carry_in[20]);
carry_in[21] = (g[20]|carry_in[20]&p[20]);
carry_out[21] = (g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))));
g[21] = a[21]&b[21];
p[21] = a[21]^b[21];

sum[21]= (p[21]^carry_in[21]);
carry_in[22] = (g[21]|carry_in[21]&p[21]);
carry_out[22] = (g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))));
g[22] = a[22]&b[22];
p[22] = a[22]^b[22];

sum[22]= (p[22]^carry_in[22]);
carry_in[23] = (g[22]|carry_in[22]&p[22]);
carry_out[23] = (g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))));
g[23] = a[23]&b[23];
p[23] = a[23]^b[23];

sum[23]= (p[23]^carry_in[23]);
carry_in[24] = (g[23]|carry_in[23]&p[23]);
carry_out[24] = (g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))));
g[24] = a[24]&b[24];
p[24] = a[24]^b[24];

sum[24]= (p[24]^carry_in[24]);
carry_in[25] = (g[24]|carry_in[24]&p[24]);
carry_out[25] = (g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))));
g[25] = a[25]&b[25];
p[25] = a[25]^b[25];

sum[25]= (p[25]^carry_in[25]);
carry_in[26] = (g[25]|carry_in[25]&p[25]);
carry_out[26] = (g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))));
g[26] = a[26]&b[26];
p[26] = a[26]^b[26];

sum[26]= (p[26]^carry_in[26]);
carry_in[27] = (g[26]|carry_in[26]&p[26]);
carry_out[27] = (g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))));
g[27] = a[27]&b[27];
p[27] = a[27]^b[27];

sum[27]= (p[27]^carry_in[27]);
carry_in[28] = (g[27]|carry_in[27]&p[27]);
carry_out[28] = (g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))));
g[28] = a[28]&b[28];
p[28] = a[28]^b[28];

sum[28]= (p[28]^carry_in[28]);
carry_in[29] = (g[28]|carry_in[28]&p[28]);
carry_out[29] = (g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))));
g[29] = a[29]&b[29];
p[29] = a[29]^b[29];

sum[29]= (p[29]^carry_in[29]);
carry_in[30] = (g[29]|carry_in[29]&p[29]);
carry_out[30] = (g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))));
g[30] = a[30]&b[30];
p[30] = a[30]^b[30];

sum[30]= (p[30]^carry_in[30]);
carry_in[31] = (g[30]|carry_in[30]&p[30]);
carry_out[31] = (g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))));
g[31] = a[31]&b[31];
p[31] = a[31]^b[31];

sum[31]= (p[31]^carry_in[31]);
carry_in[32] = (g[31]|carry_in[31]&p[31]);
carry_out[32] = (g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))));
g[32] = a[32]&b[32];
p[32] = a[32]^b[32];

sum[32]= (p[32]^carry_in[32]);
carry_in[33] = (g[32]|carry_in[32]&p[32]);
carry_out[33] = (g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))));
g[33] = a[33]&b[33];
p[33] = a[33]^b[33];

sum[33]= (p[33]^carry_in[33]);
carry_in[34] = (g[33]|carry_in[33]&p[33]);
carry_out[34] = (g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))));
g[34] = a[34]&b[34];
p[34] = a[34]^b[34];

sum[34]= (p[34]^carry_in[34]);
carry_in[35] = (g[34]|carry_in[34]&p[34]);
carry_out[35] = (g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))));
g[35] = a[35]&b[35];
p[35] = a[35]^b[35];

sum[35]= (p[35]^carry_in[35]);
carry_in[36] = (g[35]|carry_in[35]&p[35]);
carry_out[36] = (g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))));
g[36] = a[36]&b[36];
p[36] = a[36]^b[36];

sum[36]= (p[36]^carry_in[36]);
carry_in[37] = (g[36]|carry_in[36]&p[36]);
carry_out[37] = (g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))));
g[37] = a[37]&b[37];
p[37] = a[37]^b[37];

sum[37]= (p[37]^carry_in[37]);
carry_in[38] = (g[37]|carry_in[37]&p[37]);
carry_out[38] = (g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))));
g[38] = a[38]&b[38];
p[38] = a[38]^b[38];

sum[38]= (p[38]^carry_in[38]);
carry_in[39] = (g[38]|carry_in[38]&p[38]);
carry_out[39] = (g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))));
g[39] = a[39]&b[39];
p[39] = a[39]^b[39];

sum[39]= (p[39]^carry_in[39]);
carry_in[40] = (g[39]|carry_in[39]&p[39]);
carry_out[40] = (g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))));
g[40] = a[40]&b[40];
p[40] = a[40]^b[40];

sum[40]= (p[40]^carry_in[40]);
carry_in[41] = (g[40]|carry_in[40]&p[40]);
carry_out[41] = (g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))));
g[41] = a[41]&b[41];
p[41] = a[41]^b[41];

sum[41]= (p[41]^carry_in[41]);
carry_in[42] = (g[41]|carry_in[41]&p[41]);
carry_out[42] = (g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))));
g[42] = a[42]&b[42];
p[42] = a[42]^b[42];

sum[42]= (p[42]^carry_in[42]);
carry_in[43] = (g[42]|carry_in[42]&p[42]);
carry_out[43] = (g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))));
g[43] = a[43]&b[43];
p[43] = a[43]^b[43];

sum[43]= (p[43]^carry_in[43]);
carry_in[44] = (g[43]|carry_in[43]&p[43]);
carry_out[44] = (g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))));
g[44] = a[44]&b[44];
p[44] = a[44]^b[44];

sum[44]= (p[44]^carry_in[44]);
carry_in[45] = (g[44]|carry_in[44]&p[44]);
carry_out[45] = (g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))));
g[45] = a[45]&b[45];
p[45] = a[45]^b[45];

sum[45]= (p[45]^carry_in[45]);
carry_in[46] = (g[45]|carry_in[45]&p[45]);
carry_out[46] = (g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))));
g[46] = a[46]&b[46];
p[46] = a[46]^b[46];

sum[46]= (p[46]^carry_in[46]);
carry_in[47] = (g[46]|carry_in[46]&p[46]);
carry_out[47] = (g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))));
g[47] = a[47]&b[47];
p[47] = a[47]^b[47];

sum[47]= (p[47]^carry_in[47]);
carry_in[48] = (g[47]|carry_in[47]&p[47]);
carry_out[48] = (g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))));
g[48] = a[48]&b[48];
p[48] = a[48]^b[48];

sum[48]= (p[48]^carry_in[48]);
carry_in[49] = (g[48]|carry_in[48]&p[48]);
carry_out[49] = (g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))));
g[49] = a[49]&b[49];
p[49] = a[49]^b[49];

sum[49]= (p[49]^carry_in[49]);
carry_in[50] = (g[49]|carry_in[49]&p[49]);
carry_out[50] = (g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))));
g[50] = a[50]&b[50];
p[50] = a[50]^b[50];

sum[50]= (p[50]^carry_in[50]);
carry_in[51] = (g[50]|carry_in[50]&p[50]);
carry_out[51] = (g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))));
g[51] = a[51]&b[51];
p[51] = a[51]^b[51];

sum[51]= (p[51]^carry_in[51]);
carry_in[52] = (g[51]|carry_in[51]&p[51]);
carry_out[52] = (g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))));
g[52] = a[52]&b[52];
p[52] = a[52]^b[52];

sum[52]= (p[52]^carry_in[52]);
carry_in[53] = (g[52]|carry_in[52]&p[52]);
carry_out[53] = (g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))));
g[53] = a[53]&b[53];
p[53] = a[53]^b[53];

sum[53]= (p[53]^carry_in[53]);
carry_in[54] = (g[53]|carry_in[53]&p[53]);
carry_out[54] = (g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[54] = a[54]&b[54];
p[54] = a[54]^b[54];

sum[54]= (p[54]^carry_in[54]);
carry_in[55] = (g[54]|carry_in[54]&p[54]);
carry_out[55] = (g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[55] = a[55]&b[55];
p[55] = a[55]^b[55];

sum[55]= (p[55]^carry_in[55]);
carry_in[56] = (g[55]|carry_in[55]&p[55]);
carry_out[56] = (g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[56] = a[56]&b[56];
p[56] = a[56]^b[56];

sum[56]= (p[56]^carry_in[56]);
carry_in[57] = (g[56]|carry_in[56]&p[56]);
carry_out[57] = (g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[57] = a[57]&b[57];
p[57] = a[57]^b[57];

sum[57]= (p[57]^carry_in[57]);
carry_in[58] = (g[57]|carry_in[57]&p[57]);
carry_out[58] = (g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[58] = a[58]&b[58];
p[58] = a[58]^b[58];

sum[58]= (p[58]^carry_in[58]);
carry_in[59] = (g[58]|carry_in[58]&p[58]);
carry_out[59] = (g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[59] = a[59]&b[59];
p[59] = a[59]^b[59];

sum[59]= (p[59]^carry_in[59]);
carry_in[60] = (g[59]|carry_in[59]&p[59]);
carry_out[60] = (g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[60] = a[60]&b[60];
p[60] = a[60]^b[60];

sum[60]= (p[60]^carry_in[60]);
carry_in[61] = (g[60]|carry_in[60]&p[60]);
carry_out[61] = (g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[61] = a[61]&b[61];
p[61] = a[61]^b[61];

sum[61]= (p[61]^carry_in[61]);
carry_in[62] = (g[61]|carry_in[61]&p[61]);
carry_out[62] = (g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[62] = a[62]&b[62];
p[62] = a[62]^b[62];

sum[62]= (p[62]^carry_in[62]);
carry_in[63] = (g[62]|carry_in[62]&p[62]);
carry_out[63] = (g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[63] = a[63]&b[63];
p[63] = a[63]^b[63];

sum[63]= (p[63]^carry_in[63]);
carry_in[64] = (g[63]|carry_in[63]&p[63]);
carry_out[64] = (g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[64] = a[64]&b[64];
p[64] = a[64]^b[64];

sum[64]= (p[64]^carry_in[64]);
carry_in[65] = (g[64]|carry_in[64]&p[64]);
carry_out[65] = (g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[65] = a[65]&b[65];
p[65] = a[65]^b[65];

sum[65]= (p[65]^carry_in[65]);
carry_in[66] = (g[65]|carry_in[65]&p[65]);
carry_out[66] = (g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[66] = a[66]&b[66];
p[66] = a[66]^b[66];

sum[66]= (p[66]^carry_in[66]);
carry_in[67] = (g[66]|carry_in[66]&p[66]);
carry_out[67] = (g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[67] = a[67]&b[67];
p[67] = a[67]^b[67];

sum[67]= (p[67]^carry_in[67]);
carry_in[68] = (g[67]|carry_in[67]&p[67]);
carry_out[68] = (g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[68] = a[68]&b[68];
p[68] = a[68]^b[68];

sum[68]= (p[68]^carry_in[68]);
carry_in[69] = (g[68]|carry_in[68]&p[68]);
carry_out[69] = (g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[69] = a[69]&b[69];
p[69] = a[69]^b[69];

sum[69]= (p[69]^carry_in[69]);
carry_in[70] = (g[69]|carry_in[69]&p[69]);
carry_out[70] = (g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[70] = a[70]&b[70];
p[70] = a[70]^b[70];

sum[70]= (p[70]^carry_in[70]);
carry_in[71] = (g[70]|carry_in[70]&p[70]);
carry_out[71] = (g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[71] = a[71]&b[71];
p[71] = a[71]^b[71];

sum[71]= (p[71]^carry_in[71]);
carry_in[72] = (g[71]|carry_in[71]&p[71]);
carry_out[72] = (g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[72] = a[72]&b[72];
p[72] = a[72]^b[72];

sum[72]= (p[72]^carry_in[72]);
carry_in[73] = (g[72]|carry_in[72]&p[72]);
carry_out[73] = (g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[73] = a[73]&b[73];
p[73] = a[73]^b[73];

sum[73]= (p[73]^carry_in[73]);
carry_in[74] = (g[73]|carry_in[73]&p[73]);
carry_out[74] = (g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[74] = a[74]&b[74];
p[74] = a[74]^b[74];

sum[74]= (p[74]^carry_in[74]);
carry_in[75] = (g[74]|carry_in[74]&p[74]);
carry_out[75] = (g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[75] = a[75]&b[75];
p[75] = a[75]^b[75];

sum[75]= (p[75]^carry_in[75]);
carry_in[76] = (g[75]|carry_in[75]&p[75]);
carry_out[76] = (g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[76] = a[76]&b[76];
p[76] = a[76]^b[76];

sum[76]= (p[76]^carry_in[76]);
carry_in[77] = (g[76]|carry_in[76]&p[76]);
carry_out[77] = (g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[77] = a[77]&b[77];
p[77] = a[77]^b[77];

sum[77]= (p[77]^carry_in[77]);
carry_in[78] = (g[77]|carry_in[77]&p[77]);
carry_out[78] = (g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[78] = a[78]&b[78];
p[78] = a[78]^b[78];

sum[78]= (p[78]^carry_in[78]);
carry_in[79] = (g[78]|carry_in[78]&p[78]);
carry_out[79] = (g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[79] = a[79]&b[79];
p[79] = a[79]^b[79];

sum[79]= (p[79]^carry_in[79]);
carry_in[80] = (g[79]|carry_in[79]&p[79]);
carry_out[80] = (g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[80] = a[80]&b[80];
p[80] = a[80]^b[80];

sum[80]= (p[80]^carry_in[80]);
carry_in[81] = (g[80]|carry_in[80]&p[80]);
carry_out[81] = (g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[81] = a[81]&b[81];
p[81] = a[81]^b[81];

sum[81]= (p[81]^carry_in[81]);
carry_in[82] = (g[81]|carry_in[81]&p[81]);
carry_out[82] = (g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[82] = a[82]&b[82];
p[82] = a[82]^b[82];

sum[82]= (p[82]^carry_in[82]);
carry_in[83] = (g[82]|carry_in[82]&p[82]);
carry_out[83] = (g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[83] = a[83]&b[83];
p[83] = a[83]^b[83];

sum[83]= (p[83]^carry_in[83]);
carry_in[84] = (g[83]|carry_in[83]&p[83]);
carry_out[84] = (g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[84] = a[84]&b[84];
p[84] = a[84]^b[84];

sum[84]= (p[84]^carry_in[84]);
carry_in[85] = (g[84]|carry_in[84]&p[84]);
carry_out[85] = (g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[85] = a[85]&b[85];
p[85] = a[85]^b[85];

sum[85]= (p[85]^carry_in[85]);
carry_in[86] = (g[85]|carry_in[85]&p[85]);
carry_out[86] = (g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[86] = a[86]&b[86];
p[86] = a[86]^b[86];

sum[86]= (p[86]^carry_in[86]);
carry_in[87] = (g[86]|carry_in[86]&p[86]);
carry_out[87] = (g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[87] = a[87]&b[87];
p[87] = a[87]^b[87];

sum[87]= (p[87]^carry_in[87]);
carry_in[88] = (g[87]|carry_in[87]&p[87]);
carry_out[88] = (g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[88] = a[88]&b[88];
p[88] = a[88]^b[88];

sum[88]= (p[88]^carry_in[88]);
carry_in[89] = (g[88]|carry_in[88]&p[88]);
carry_out[89] = (g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[89] = a[89]&b[89];
p[89] = a[89]^b[89];

sum[89]= (p[89]^carry_in[89]);
carry_in[90] = (g[89]|carry_in[89]&p[89]);
carry_out[90] = (g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[90] = a[90]&b[90];
p[90] = a[90]^b[90];

sum[90]= (p[90]^carry_in[90]);
carry_in[91] = (g[90]|carry_in[90]&p[90]);
carry_out[91] = (g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[91] = a[91]&b[91];
p[91] = a[91]^b[91];

sum[91]= (p[91]^carry_in[91]);
carry_in[92] = (g[91]|carry_in[91]&p[91]);
carry_out[92] = (g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[92] = a[92]&b[92];
p[92] = a[92]^b[92];

sum[92]= (p[92]^carry_in[92]);
carry_in[93] = (g[92]|carry_in[92]&p[92]);
carry_out[93] = (g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[93] = a[93]&b[93];
p[93] = a[93]^b[93];

sum[93]= (p[93]^carry_in[93]);
carry_in[94] = (g[93]|carry_in[93]&p[93]);
carry_out[94] = (g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[94] = a[94]&b[94];
p[94] = a[94]^b[94];

sum[94]= (p[94]^carry_in[94]);
carry_in[95] = (g[94]|carry_in[94]&p[94]);
carry_out[95] = (g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[95] = a[95]&b[95];
p[95] = a[95]^b[95];

sum[95]= (p[95]^carry_in[95]);
carry_in[96] = (g[95]|carry_in[95]&p[95]);
carry_out[96] = (g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[96] = a[96]&b[96];
p[96] = a[96]^b[96];

sum[96]= (p[96]^carry_in[96]);
carry_in[97] = (g[96]|carry_in[96]&p[96]);
carry_out[97] = (g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[97] = a[97]&b[97];
p[97] = a[97]^b[97];

sum[97]= (p[97]^carry_in[97]);
carry_in[98] = (g[97]|carry_in[97]&p[97]);
carry_out[98] = (g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[98] = a[98]&b[98];
p[98] = a[98]^b[98];

sum[98]= (p[98]^carry_in[98]);
carry_in[99] = (g[98]|carry_in[98]&p[98]);
carry_out[99] = (g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[99] = a[99]&b[99];
p[99] = a[99]^b[99];

sum[99]= (p[99]^carry_in[99]);
carry_in[100] = (g[99]|carry_in[99]&p[99]);
carry_out[100] = (g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[100] = a[100]&b[100];
p[100] = a[100]^b[100];

sum[100]= (p[100]^carry_in[100]);
carry_in[101] = (g[100]|carry_in[100]&p[100]);
carry_out[101] = (g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[101] = a[101]&b[101];
p[101] = a[101]^b[101];

sum[101]= (p[101]^carry_in[101]);
carry_in[102] = (g[101]|carry_in[101]&p[101]);
carry_out[102] = (g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[102] = a[102]&b[102];
p[102] = a[102]^b[102];

sum[102]= (p[102]^carry_in[102]);
carry_in[103] = (g[102]|carry_in[102]&p[102]);
carry_out[103] = (g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[103] = a[103]&b[103];
p[103] = a[103]^b[103];

sum[103]= (p[103]^carry_in[103]);
carry_in[104] = (g[103]|carry_in[103]&p[103]);
carry_out[104] = (g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[104] = a[104]&b[104];
p[104] = a[104]^b[104];

sum[104]= (p[104]^carry_in[104]);
carry_in[105] = (g[104]|carry_in[104]&p[104]);
carry_out[105] = (g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[105] = a[105]&b[105];
p[105] = a[105]^b[105];

sum[105]= (p[105]^carry_in[105]);
carry_in[106] = (g[105]|carry_in[105]&p[105]);
carry_out[106] = (g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[106] = a[106]&b[106];
p[106] = a[106]^b[106];

sum[106]= (p[106]^carry_in[106]);
carry_in[107] = (g[106]|carry_in[106]&p[106]);
carry_out[107] = (g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[107] = a[107]&b[107];
p[107] = a[107]^b[107];

sum[107]= (p[107]^carry_in[107]);
carry_in[108] = (g[107]|carry_in[107]&p[107]);
carry_out[108] = (g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[108] = a[108]&b[108];
p[108] = a[108]^b[108];

sum[108]= (p[108]^carry_in[108]);
carry_in[109] = (g[108]|carry_in[108]&p[108]);
carry_out[109] = (g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[109] = a[109]&b[109];
p[109] = a[109]^b[109];

sum[109]= (p[109]^carry_in[109]);
carry_in[110] = (g[109]|carry_in[109]&p[109]);
carry_out[110] = (g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[110] = a[110]&b[110];
p[110] = a[110]^b[110];

sum[110]= (p[110]^carry_in[110]);
carry_in[111] = (g[110]|carry_in[110]&p[110]);
carry_out[111] = (g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[111] = a[111]&b[111];
p[111] = a[111]^b[111];

sum[111]= (p[111]^carry_in[111]);
carry_in[112] = (g[111]|carry_in[111]&p[111]);
carry_out[112] = (g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[112] = a[112]&b[112];
p[112] = a[112]^b[112];

sum[112]= (p[112]^carry_in[112]);
carry_in[113] = (g[112]|carry_in[112]&p[112]);
carry_out[113] = (g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[113] = a[113]&b[113];
p[113] = a[113]^b[113];

sum[113]= (p[113]^carry_in[113]);
carry_in[114] = (g[113]|carry_in[113]&p[113]);
carry_out[114] = (g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[114] = a[114]&b[114];
p[114] = a[114]^b[114];

sum[114]= (p[114]^carry_in[114]);
carry_in[115] = (g[114]|carry_in[114]&p[114]);
carry_out[115] = (g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[115] = a[115]&b[115];
p[115] = a[115]^b[115];

sum[115]= (p[115]^carry_in[115]);
carry_in[116] = (g[115]|carry_in[115]&p[115]);
carry_out[116] = (g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[116] = a[116]&b[116];
p[116] = a[116]^b[116];

sum[116]= (p[116]^carry_in[116]);
carry_in[117] = (g[116]|carry_in[116]&p[116]);
carry_out[117] = (g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[117] = a[117]&b[117];
p[117] = a[117]^b[117];

sum[117]= (p[117]^carry_in[117]);
carry_in[118] = (g[117]|carry_in[117]&p[117]);
carry_out[118] = (g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[118] = a[118]&b[118];
p[118] = a[118]^b[118];

sum[118]= (p[118]^carry_in[118]);
carry_in[119] = (g[118]|carry_in[118]&p[118]);
carry_out[119] = (g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[119] = a[119]&b[119];
p[119] = a[119]^b[119];

sum[119]= (p[119]^carry_in[119]);
carry_in[120] = (g[119]|carry_in[119]&p[119]);
carry_out[120] = (g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[120] = a[120]&b[120];
p[120] = a[120]^b[120];

sum[120]= (p[120]^carry_in[120]);
carry_in[121] = (g[120]|carry_in[120]&p[120]);
carry_out[121] = (g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[121] = a[121]&b[121];
p[121] = a[121]^b[121];

sum[121]= (p[121]^carry_in[121]);
carry_in[122] = (g[121]|carry_in[121]&p[121]);
carry_out[122] = (g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[122] = a[122]&b[122];
p[122] = a[122]^b[122];

sum[122]= (p[122]^carry_in[122]);
carry_in[123] = (g[122]|carry_in[122]&p[122]);
carry_out[123] = (g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[123] = a[123]&b[123];
p[123] = a[123]^b[123];

sum[123]= (p[123]^carry_in[123]);
carry_in[124] = (g[123]|carry_in[123]&p[123]);
carry_out[124] = (g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[124] = a[124]&b[124];
p[124] = a[124]^b[124];

sum[124]= (p[124]^carry_in[124]);
carry_in[125] = (g[124]|carry_in[124]&p[124]);
carry_out[125] = (g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[125] = a[125]&b[125];
p[125] = a[125]^b[125];

sum[125]= (p[125]^carry_in[125]);
carry_in[126] = (g[125]|carry_in[125]&p[125]);
carry_out[126] = (g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[126] = a[126]&b[126];
p[126] = a[126]^b[126];

sum[126]= (p[126]^carry_in[126]);
carry_in[127] = (g[126]|carry_in[126]&p[126]);
carry_out[127] = (g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[127] = a[127]&b[127];
p[127] = a[127]^b[127];

sum[127]= (p[127]^carry_in[127]);
carry_in[128] = (g[127]|carry_in[127]&p[127]);
carry_out[128] = (g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[128] = a[128]&b[128];
p[128] = a[128]^b[128];

sum[128]= (p[128]^carry_in[128]);
carry_in[129] = (g[128]|carry_in[128]&p[128]);
carry_out[129] = (g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[129] = a[129]&b[129];
p[129] = a[129]^b[129];

sum[129]= (p[129]^carry_in[129]);
carry_in[130] = (g[129]|carry_in[129]&p[129]);
carry_out[130] = (g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[130] = a[130]&b[130];
p[130] = a[130]^b[130];

sum[130]= (p[130]^carry_in[130]);
carry_in[131] = (g[130]|carry_in[130]&p[130]);
carry_out[131] = (g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[131] = a[131]&b[131];
p[131] = a[131]^b[131];

sum[131]= (p[131]^carry_in[131]);
carry_in[132] = (g[131]|carry_in[131]&p[131]);
carry_out[132] = (g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[132] = a[132]&b[132];
p[132] = a[132]^b[132];

sum[132]= (p[132]^carry_in[132]);
carry_in[133] = (g[132]|carry_in[132]&p[132]);
carry_out[133] = (g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[133] = a[133]&b[133];
p[133] = a[133]^b[133];

sum[133]= (p[133]^carry_in[133]);
carry_in[134] = (g[133]|carry_in[133]&p[133]);
carry_out[134] = (g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[134] = a[134]&b[134];
p[134] = a[134]^b[134];

sum[134]= (p[134]^carry_in[134]);
carry_in[135] = (g[134]|carry_in[134]&p[134]);
carry_out[135] = (g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[135] = a[135]&b[135];
p[135] = a[135]^b[135];

sum[135]= (p[135]^carry_in[135]);
carry_in[136] = (g[135]|carry_in[135]&p[135]);
carry_out[136] = (g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[136] = a[136]&b[136];
p[136] = a[136]^b[136];

sum[136]= (p[136]^carry_in[136]);
carry_in[137] = (g[136]|carry_in[136]&p[136]);
carry_out[137] = (g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[137] = a[137]&b[137];
p[137] = a[137]^b[137];

sum[137]= (p[137]^carry_in[137]);
carry_in[138] = (g[137]|carry_in[137]&p[137]);
carry_out[138] = (g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[138] = a[138]&b[138];
p[138] = a[138]^b[138];

sum[138]= (p[138]^carry_in[138]);
carry_in[139] = (g[138]|carry_in[138]&p[138]);
carry_out[139] = (g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[139] = a[139]&b[139];
p[139] = a[139]^b[139];

sum[139]= (p[139]^carry_in[139]);
carry_in[140] = (g[139]|carry_in[139]&p[139]);
carry_out[140] = (g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[140] = a[140]&b[140];
p[140] = a[140]^b[140];

sum[140]= (p[140]^carry_in[140]);
carry_in[141] = (g[140]|carry_in[140]&p[140]);
carry_out[141] = (g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[141] = a[141]&b[141];
p[141] = a[141]^b[141];

sum[141]= (p[141]^carry_in[141]);
carry_in[142] = (g[141]|carry_in[141]&p[141]);
carry_out[142] = (g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[142] = a[142]&b[142];
p[142] = a[142]^b[142];

sum[142]= (p[142]^carry_in[142]);
carry_in[143] = (g[142]|carry_in[142]&p[142]);
carry_out[143] = (g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[143] = a[143]&b[143];
p[143] = a[143]^b[143];

sum[143]= (p[143]^carry_in[143]);
carry_in[144] = (g[143]|carry_in[143]&p[143]);
carry_out[144] = (g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[144] = a[144]&b[144];
p[144] = a[144]^b[144];

sum[144]= (p[144]^carry_in[144]);
carry_in[145] = (g[144]|carry_in[144]&p[144]);
carry_out[145] = (g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[145] = a[145]&b[145];
p[145] = a[145]^b[145];

sum[145]= (p[145]^carry_in[145]);
carry_in[146] = (g[145]|carry_in[145]&p[145]);
carry_out[146] = (g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[146] = a[146]&b[146];
p[146] = a[146]^b[146];

sum[146]= (p[146]^carry_in[146]);
carry_in[147] = (g[146]|carry_in[146]&p[146]);
carry_out[147] = (g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[147] = a[147]&b[147];
p[147] = a[147]^b[147];

sum[147]= (p[147]^carry_in[147]);
carry_in[148] = (g[147]|carry_in[147]&p[147]);
carry_out[148] = (g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[148] = a[148]&b[148];
p[148] = a[148]^b[148];

sum[148]= (p[148]^carry_in[148]);
carry_in[149] = (g[148]|carry_in[148]&p[148]);
carry_out[149] = (g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[149] = a[149]&b[149];
p[149] = a[149]^b[149];

sum[149]= (p[149]^carry_in[149]);
carry_in[150] = (g[149]|carry_in[149]&p[149]);
carry_out[150] = (g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[150] = a[150]&b[150];
p[150] = a[150]^b[150];

sum[150]= (p[150]^carry_in[150]);
carry_in[151] = (g[150]|carry_in[150]&p[150]);
carry_out[151] = (g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[151] = a[151]&b[151];
p[151] = a[151]^b[151];

sum[151]= (p[151]^carry_in[151]);
carry_in[152] = (g[151]|carry_in[151]&p[151]);
carry_out[152] = (g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[152] = a[152]&b[152];
p[152] = a[152]^b[152];

sum[152]= (p[152]^carry_in[152]);
carry_in[153] = (g[152]|carry_in[152]&p[152]);
carry_out[153] = (g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[153] = a[153]&b[153];
p[153] = a[153]^b[153];

sum[153]= (p[153]^carry_in[153]);
carry_in[154] = (g[153]|carry_in[153]&p[153]);
carry_out[154] = (g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[154] = a[154]&b[154];
p[154] = a[154]^b[154];

sum[154]= (p[154]^carry_in[154]);
carry_in[155] = (g[154]|carry_in[154]&p[154]);
carry_out[155] = (g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[155] = a[155]&b[155];
p[155] = a[155]^b[155];

sum[155]= (p[155]^carry_in[155]);
carry_in[156] = (g[155]|carry_in[155]&p[155]);
carry_out[156] = (g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[156] = a[156]&b[156];
p[156] = a[156]^b[156];

sum[156]= (p[156]^carry_in[156]);
carry_in[157] = (g[156]|carry_in[156]&p[156]);
carry_out[157] = (g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[157] = a[157]&b[157];
p[157] = a[157]^b[157];

sum[157]= (p[157]^carry_in[157]);
carry_in[158] = (g[157]|carry_in[157]&p[157]);
carry_out[158] = (g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[158] = a[158]&b[158];
p[158] = a[158]^b[158];

sum[158]= (p[158]^carry_in[158]);
carry_in[159] = (g[158]|carry_in[158]&p[158]);
carry_out[159] = (g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[159] = a[159]&b[159];
p[159] = a[159]^b[159];

sum[159]= (p[159]^carry_in[159]);
carry_in[160] = (g[159]|carry_in[159]&p[159]);
carry_out[160] = (g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[160] = a[160]&b[160];
p[160] = a[160]^b[160];

sum[160]= (p[160]^carry_in[160]);
carry_in[161] = (g[160]|carry_in[160]&p[160]);
carry_out[161] = (g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[161] = a[161]&b[161];
p[161] = a[161]^b[161];

sum[161]= (p[161]^carry_in[161]);
carry_in[162] = (g[161]|carry_in[161]&p[161]);
carry_out[162] = (g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[162] = a[162]&b[162];
p[162] = a[162]^b[162];

sum[162]= (p[162]^carry_in[162]);
carry_in[163] = (g[162]|carry_in[162]&p[162]);
carry_out[163] = (g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[163] = a[163]&b[163];
p[163] = a[163]^b[163];

sum[163]= (p[163]^carry_in[163]);
carry_in[164] = (g[163]|carry_in[163]&p[163]);
carry_out[164] = (g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[164] = a[164]&b[164];
p[164] = a[164]^b[164];

sum[164]= (p[164]^carry_in[164]);
carry_in[165] = (g[164]|carry_in[164]&p[164]);
carry_out[165] = (g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[165] = a[165]&b[165];
p[165] = a[165]^b[165];

sum[165]= (p[165]^carry_in[165]);
carry_in[166] = (g[165]|carry_in[165]&p[165]);
carry_out[166] = (g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[166] = a[166]&b[166];
p[166] = a[166]^b[166];

sum[166]= (p[166]^carry_in[166]);
carry_in[167] = (g[166]|carry_in[166]&p[166]);
carry_out[167] = (g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[167] = a[167]&b[167];
p[167] = a[167]^b[167];

sum[167]= (p[167]^carry_in[167]);
carry_in[168] = (g[167]|carry_in[167]&p[167]);
carry_out[168] = (g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[168] = a[168]&b[168];
p[168] = a[168]^b[168];

sum[168]= (p[168]^carry_in[168]);
carry_in[169] = (g[168]|carry_in[168]&p[168]);
carry_out[169] = (g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[169] = a[169]&b[169];
p[169] = a[169]^b[169];

sum[169]= (p[169]^carry_in[169]);
carry_in[170] = (g[169]|carry_in[169]&p[169]);
carry_out[170] = (g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[170] = a[170]&b[170];
p[170] = a[170]^b[170];

sum[170]= (p[170]^carry_in[170]);
carry_in[171] = (g[170]|carry_in[170]&p[170]);
carry_out[171] = (g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[171] = a[171]&b[171];
p[171] = a[171]^b[171];

sum[171]= (p[171]^carry_in[171]);
carry_in[172] = (g[171]|carry_in[171]&p[171]);
carry_out[172] = (g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[172] = a[172]&b[172];
p[172] = a[172]^b[172];

sum[172]= (p[172]^carry_in[172]);
carry_in[173] = (g[172]|carry_in[172]&p[172]);
carry_out[173] = (g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[173] = a[173]&b[173];
p[173] = a[173]^b[173];

sum[173]= (p[173]^carry_in[173]);
carry_in[174] = (g[173]|carry_in[173]&p[173]);
carry_out[174] = (g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[174] = a[174]&b[174];
p[174] = a[174]^b[174];

sum[174]= (p[174]^carry_in[174]);
carry_in[175] = (g[174]|carry_in[174]&p[174]);
carry_out[175] = (g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[175] = a[175]&b[175];
p[175] = a[175]^b[175];

sum[175]= (p[175]^carry_in[175]);
carry_in[176] = (g[175]|carry_in[175]&p[175]);
carry_out[176] = (g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[176] = a[176]&b[176];
p[176] = a[176]^b[176];

sum[176]= (p[176]^carry_in[176]);
carry_in[177] = (g[176]|carry_in[176]&p[176]);
carry_out[177] = (g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[177] = a[177]&b[177];
p[177] = a[177]^b[177];

sum[177]= (p[177]^carry_in[177]);
carry_in[178] = (g[177]|carry_in[177]&p[177]);
carry_out[178] = (g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[178] = a[178]&b[178];
p[178] = a[178]^b[178];

sum[178]= (p[178]^carry_in[178]);
carry_in[179] = (g[178]|carry_in[178]&p[178]);
carry_out[179] = (g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[179] = a[179]&b[179];
p[179] = a[179]^b[179];

sum[179]= (p[179]^carry_in[179]);
carry_in[180] = (g[179]|carry_in[179]&p[179]);
carry_out[180] = (g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[180] = a[180]&b[180];
p[180] = a[180]^b[180];

sum[180]= (p[180]^carry_in[180]);
carry_in[181] = (g[180]|carry_in[180]&p[180]);
carry_out[181] = (g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[181] = a[181]&b[181];
p[181] = a[181]^b[181];

sum[181]= (p[181]^carry_in[181]);
carry_in[182] = (g[181]|carry_in[181]&p[181]);
carry_out[182] = (g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[182] = a[182]&b[182];
p[182] = a[182]^b[182];

sum[182]= (p[182]^carry_in[182]);
carry_in[183] = (g[182]|carry_in[182]&p[182]);
carry_out[183] = (g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[183] = a[183]&b[183];
p[183] = a[183]^b[183];

sum[183]= (p[183]^carry_in[183]);
carry_in[184] = (g[183]|carry_in[183]&p[183]);
carry_out[184] = (g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[184] = a[184]&b[184];
p[184] = a[184]^b[184];

sum[184]= (p[184]^carry_in[184]);
carry_in[185] = (g[184]|carry_in[184]&p[184]);
carry_out[185] = (g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[185] = a[185]&b[185];
p[185] = a[185]^b[185];

sum[185]= (p[185]^carry_in[185]);
carry_in[186] = (g[185]|carry_in[185]&p[185]);
carry_out[186] = (g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[186] = a[186]&b[186];
p[186] = a[186]^b[186];

sum[186]= (p[186]^carry_in[186]);
carry_in[187] = (g[186]|carry_in[186]&p[186]);
carry_out[187] = (g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[187] = a[187]&b[187];
p[187] = a[187]^b[187];

sum[187]= (p[187]^carry_in[187]);
carry_in[188] = (g[187]|carry_in[187]&p[187]);
carry_out[188] = (g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[188] = a[188]&b[188];
p[188] = a[188]^b[188];

sum[188]= (p[188]^carry_in[188]);
carry_in[189] = (g[188]|carry_in[188]&p[188]);
carry_out[189] = (g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[189] = a[189]&b[189];
p[189] = a[189]^b[189];

sum[189]= (p[189]^carry_in[189]);
carry_in[190] = (g[189]|carry_in[189]&p[189]);
carry_out[190] = (g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[190] = a[190]&b[190];
p[190] = a[190]^b[190];

sum[190]= (p[190]^carry_in[190]);
carry_in[191] = (g[190]|carry_in[190]&p[190]);
carry_out[191] = (g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[191] = a[191]&b[191];
p[191] = a[191]^b[191];

sum[191]= (p[191]^carry_in[191]);
carry_in[192] = (g[191]|carry_in[191]&p[191]);
carry_out[192] = (g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[192] = a[192]&b[192];
p[192] = a[192]^b[192];

sum[192]= (p[192]^carry_in[192]);
carry_in[193] = (g[192]|carry_in[192]&p[192]);
carry_out[193] = (g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[193] = a[193]&b[193];
p[193] = a[193]^b[193];

sum[193]= (p[193]^carry_in[193]);
carry_in[194] = (g[193]|carry_in[193]&p[193]);
carry_out[194] = (g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[194] = a[194]&b[194];
p[194] = a[194]^b[194];

sum[194]= (p[194]^carry_in[194]);
carry_in[195] = (g[194]|carry_in[194]&p[194]);
carry_out[195] = (g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[195] = a[195]&b[195];
p[195] = a[195]^b[195];

sum[195]= (p[195]^carry_in[195]);
carry_in[196] = (g[195]|carry_in[195]&p[195]);
carry_out[196] = (g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[196] = a[196]&b[196];
p[196] = a[196]^b[196];

sum[196]= (p[196]^carry_in[196]);
carry_in[197] = (g[196]|carry_in[196]&p[196]);
carry_out[197] = (g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[197] = a[197]&b[197];
p[197] = a[197]^b[197];

sum[197]= (p[197]^carry_in[197]);
carry_in[198] = (g[197]|carry_in[197]&p[197]);
carry_out[198] = (g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[198] = a[198]&b[198];
p[198] = a[198]^b[198];

sum[198]= (p[198]^carry_in[198]);
carry_in[199] = (g[198]|carry_in[198]&p[198]);
carry_out[199] = (g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[199] = a[199]&b[199];
p[199] = a[199]^b[199];

sum[199]= (p[199]^carry_in[199]);
carry_in[200] = (g[199]|carry_in[199]&p[199]);
carry_out[200] = (g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[200] = a[200]&b[200];
p[200] = a[200]^b[200];

sum[200]= (p[200]^carry_in[200]);
carry_in[201] = (g[200]|carry_in[200]&p[200]);
carry_out[201] = (g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[201] = a[201]&b[201];
p[201] = a[201]^b[201];

sum[201]= (p[201]^carry_in[201]);
carry_in[202] = (g[201]|carry_in[201]&p[201]);
carry_out[202] = (g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[202] = a[202]&b[202];
p[202] = a[202]^b[202];

sum[202]= (p[202]^carry_in[202]);
carry_in[203] = (g[202]|carry_in[202]&p[202]);
carry_out[203] = (g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[203] = a[203]&b[203];
p[203] = a[203]^b[203];

sum[203]= (p[203]^carry_in[203]);
carry_in[204] = (g[203]|carry_in[203]&p[203]);
carry_out[204] = (g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[204] = a[204]&b[204];
p[204] = a[204]^b[204];

sum[204]= (p[204]^carry_in[204]);
carry_in[205] = (g[204]|carry_in[204]&p[204]);
carry_out[205] = (g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[205] = a[205]&b[205];
p[205] = a[205]^b[205];

sum[205]= (p[205]^carry_in[205]);
carry_in[206] = (g[205]|carry_in[205]&p[205]);
carry_out[206] = (g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[206] = a[206]&b[206];
p[206] = a[206]^b[206];

sum[206]= (p[206]^carry_in[206]);
carry_in[207] = (g[206]|carry_in[206]&p[206]);
carry_out[207] = (g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[207] = a[207]&b[207];
p[207] = a[207]^b[207];

sum[207]= (p[207]^carry_in[207]);
carry_in[208] = (g[207]|carry_in[207]&p[207]);
carry_out[208] = (g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[208] = a[208]&b[208];
p[208] = a[208]^b[208];

sum[208]= (p[208]^carry_in[208]);
carry_in[209] = (g[208]|carry_in[208]&p[208]);
carry_out[209] = (g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[209] = a[209]&b[209];
p[209] = a[209]^b[209];

sum[209]= (p[209]^carry_in[209]);
carry_in[210] = (g[209]|carry_in[209]&p[209]);
carry_out[210] = (g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[210] = a[210]&b[210];
p[210] = a[210]^b[210];

sum[210]= (p[210]^carry_in[210]);
carry_in[211] = (g[210]|carry_in[210]&p[210]);
carry_out[211] = (g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[211] = a[211]&b[211];
p[211] = a[211]^b[211];

sum[211]= (p[211]^carry_in[211]);
carry_in[212] = (g[211]|carry_in[211]&p[211]);
carry_out[212] = (g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[212] = a[212]&b[212];
p[212] = a[212]^b[212];

sum[212]= (p[212]^carry_in[212]);
carry_in[213] = (g[212]|carry_in[212]&p[212]);
carry_out[213] = (g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[213] = a[213]&b[213];
p[213] = a[213]^b[213];

sum[213]= (p[213]^carry_in[213]);
carry_in[214] = (g[213]|carry_in[213]&p[213]);
carry_out[214] = (g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[214] = a[214]&b[214];
p[214] = a[214]^b[214];

sum[214]= (p[214]^carry_in[214]);
carry_in[215] = (g[214]|carry_in[214]&p[214]);
carry_out[215] = (g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[215] = a[215]&b[215];
p[215] = a[215]^b[215];

sum[215]= (p[215]^carry_in[215]);
carry_in[216] = (g[215]|carry_in[215]&p[215]);
carry_out[216] = (g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[216] = a[216]&b[216];
p[216] = a[216]^b[216];

sum[216]= (p[216]^carry_in[216]);
carry_in[217] = (g[216]|carry_in[216]&p[216]);
carry_out[217] = (g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[217] = a[217]&b[217];
p[217] = a[217]^b[217];

sum[217]= (p[217]^carry_in[217]);
carry_in[218] = (g[217]|carry_in[217]&p[217]);
carry_out[218] = (g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[218] = a[218]&b[218];
p[218] = a[218]^b[218];

sum[218]= (p[218]^carry_in[218]);
carry_in[219] = (g[218]|carry_in[218]&p[218]);
carry_out[219] = (g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[219] = a[219]&b[219];
p[219] = a[219]^b[219];

sum[219]= (p[219]^carry_in[219]);
carry_in[220] = (g[219]|carry_in[219]&p[219]);
carry_out[220] = (g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[220] = a[220]&b[220];
p[220] = a[220]^b[220];

sum[220]= (p[220]^carry_in[220]);
carry_in[221] = (g[220]|carry_in[220]&p[220]);
carry_out[221] = (g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[221] = a[221]&b[221];
p[221] = a[221]^b[221];

sum[221]= (p[221]^carry_in[221]);
carry_in[222] = (g[221]|carry_in[221]&p[221]);
carry_out[222] = (g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[222] = a[222]&b[222];
p[222] = a[222]^b[222];

sum[222]= (p[222]^carry_in[222]);
carry_in[223] = (g[222]|carry_in[222]&p[222]);
carry_out[223] = (g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[223] = a[223]&b[223];
p[223] = a[223]^b[223];

sum[223]= (p[223]^carry_in[223]);
carry_in[224] = (g[223]|carry_in[223]&p[223]);
carry_out[224] = (g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[224] = a[224]&b[224];
p[224] = a[224]^b[224];

sum[224]= (p[224]^carry_in[224]);
carry_in[225] = (g[224]|carry_in[224]&p[224]);
carry_out[225] = (g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[225] = a[225]&b[225];
p[225] = a[225]^b[225];

sum[225]= (p[225]^carry_in[225]);
carry_in[226] = (g[225]|carry_in[225]&p[225]);
carry_out[226] = (g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[226] = a[226]&b[226];
p[226] = a[226]^b[226];

sum[226]= (p[226]^carry_in[226]);
carry_in[227] = (g[226]|carry_in[226]&p[226]);
carry_out[227] = (g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[227] = a[227]&b[227];
p[227] = a[227]^b[227];

sum[227]= (p[227]^carry_in[227]);
carry_in[228] = (g[227]|carry_in[227]&p[227]);
carry_out[228] = (g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[228] = a[228]&b[228];
p[228] = a[228]^b[228];

sum[228]= (p[228]^carry_in[228]);
carry_in[229] = (g[228]|carry_in[228]&p[228]);
carry_out[229] = (g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[229] = a[229]&b[229];
p[229] = a[229]^b[229];

sum[229]= (p[229]^carry_in[229]);
carry_in[230] = (g[229]|carry_in[229]&p[229]);
carry_out[230] = (g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[230] = a[230]&b[230];
p[230] = a[230]^b[230];

sum[230]= (p[230]^carry_in[230]);
carry_in[231] = (g[230]|carry_in[230]&p[230]);
carry_out[231] = (g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[231] = a[231]&b[231];
p[231] = a[231]^b[231];

sum[231]= (p[231]^carry_in[231]);
carry_in[232] = (g[231]|carry_in[231]&p[231]);
carry_out[232] = (g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[232] = a[232]&b[232];
p[232] = a[232]^b[232];

sum[232]= (p[232]^carry_in[232]);
carry_in[233] = (g[232]|carry_in[232]&p[232]);
carry_out[233] = (g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[233] = a[233]&b[233];
p[233] = a[233]^b[233];

sum[233]= (p[233]^carry_in[233]);
carry_in[234] = (g[233]|carry_in[233]&p[233]);
carry_out[234] = (g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[234] = a[234]&b[234];
p[234] = a[234]^b[234];

sum[234]= (p[234]^carry_in[234]);
carry_in[235] = (g[234]|carry_in[234]&p[234]);
carry_out[235] = (g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[235] = a[235]&b[235];
p[235] = a[235]^b[235];

sum[235]= (p[235]^carry_in[235]);
carry_in[236] = (g[235]|carry_in[235]&p[235]);
carry_out[236] = (g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[236] = a[236]&b[236];
p[236] = a[236]^b[236];

sum[236]= (p[236]^carry_in[236]);
carry_in[237] = (g[236]|carry_in[236]&p[236]);
carry_out[237] = (g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[237] = a[237]&b[237];
p[237] = a[237]^b[237];

sum[237]= (p[237]^carry_in[237]);
carry_in[238] = (g[237]|carry_in[237]&p[237]);
carry_out[238] = (g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[238] = a[238]&b[238];
p[238] = a[238]^b[238];

sum[238]= (p[238]^carry_in[238]);
carry_in[239] = (g[238]|carry_in[238]&p[238]);
carry_out[239] = (g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[239] = a[239]&b[239];
p[239] = a[239]^b[239];

sum[239]= (p[239]^carry_in[239]);
carry_in[240] = (g[239]|carry_in[239]&p[239]);
carry_out[240] = (g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[240] = a[240]&b[240];
p[240] = a[240]^b[240];

sum[240]= (p[240]^carry_in[240]);
carry_in[241] = (g[240]|carry_in[240]&p[240]);
carry_out[241] = (g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[241] = a[241]&b[241];
p[241] = a[241]^b[241];

sum[241]= (p[241]^carry_in[241]);
carry_in[242] = (g[241]|carry_in[241]&p[241]);
carry_out[242] = (g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[242] = a[242]&b[242];
p[242] = a[242]^b[242];

sum[242]= (p[242]^carry_in[242]);
carry_in[243] = (g[242]|carry_in[242]&p[242]);
carry_out[243] = (g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[243] = a[243]&b[243];
p[243] = a[243]^b[243];

sum[243]= (p[243]^carry_in[243]);
carry_in[244] = (g[243]|carry_in[243]&p[243]);
carry_out[244] = (g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[244] = a[244]&b[244];
p[244] = a[244]^b[244];

sum[244]= (p[244]^carry_in[244]);
carry_in[245] = (g[244]|carry_in[244]&p[244]);
carry_out[245] = (g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[245] = a[245]&b[245];
p[245] = a[245]^b[245];

sum[245]= (p[245]^carry_in[245]);
carry_in[246] = (g[245]|carry_in[245]&p[245]);
carry_out[246] = (g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[246] = a[246]&b[246];
p[246] = a[246]^b[246];

sum[246]= (p[246]^carry_in[246]);
carry_in[247] = (g[246]|carry_in[246]&p[246]);
carry_out[247] = (g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[247] = a[247]&b[247];
p[247] = a[247]^b[247];

sum[247]= (p[247]^carry_in[247]);
carry_in[248] = (g[247]|carry_in[247]&p[247]);
carry_out[248] = (g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[248] = a[248]&b[248];
p[248] = a[248]^b[248];

sum[248]= (p[248]^carry_in[248]);
carry_in[249] = (g[248]|carry_in[248]&p[248]);
carry_out[249] = (g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[249] = a[249]&b[249];
p[249] = a[249]^b[249];

sum[249]= (p[249]^carry_in[249]);
carry_in[250] = (g[249]|carry_in[249]&p[249]);
carry_out[250] = (g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[250] = a[250]&b[250];
p[250] = a[250]^b[250];

sum[250]= (p[250]^carry_in[250]);
carry_in[251] = (g[250]|carry_in[250]&p[250]);
carry_out[251] = (g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[251] = a[251]&b[251];
p[251] = a[251]^b[251];

sum[251]= (p[251]^carry_in[251]);
carry_in[252] = (g[251]|carry_in[251]&p[251]);
carry_out[252] = (g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[252] = a[252]&b[252];
p[252] = a[252]^b[252];

sum[252]= (p[252]^carry_in[252]);
carry_in[253] = (g[252]|carry_in[252]&p[252]);
carry_out[253] = (g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[253] = a[253]&b[253];
p[253] = a[253]^b[253];

sum[253]= (p[253]^carry_in[253]);
carry_in[254] = (g[253]|carry_in[253]&p[253]);
carry_out[254] = (g[253] | p[253] &(g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
g[254] = a[254]&b[254];
p[254] = a[254]^b[254];

sum[254]= (p[254]^carry_in[254]);
carry_in[255] = (g[254]|carry_in[254]&p[254]);
carry_out[255] = (g[254] | p[254] &(g[253] | p[253] &(g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0])))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));



sum[255]= ((a[255]^b[255])^carry_in[254]);
g[255] = a[255]&b[255];
p[255] = a[255]^b[255];
carry_out_overflow = (g[255] | p[255] & (g[254] | p[254] &(g[253] | p[253] &(g[252] | p[252] &(g[251] | p[251] &(g[250] | p[250] &(g[249] | p[249] &(g[248] | p[248] &(g[247] | p[247] &(g[246] | p[246] &(g[245] | p[245] &(g[244] | p[244] &(g[243] | p[243] &(g[242] | p[242] &(g[241] | p[241] &(g[240] | p[240] &(g[239] | p[239] &(g[238] | p[238] &(g[237] | p[237] &(g[236] | p[236] &(g[235] | p[235] &(g[234] | p[234] &(g[233] | p[233] &(g[232] | p[232] &(g[231] | p[231] &(g[230] | p[230] &(g[229] | p[229] &(g[228] | p[228] &(g[227] | p[227] &(g[226] | p[226] &(g[225] | p[225] &(g[224] | p[224] &(g[223] | p[223] &(g[222] | p[222] &(g[221] | p[221] &(g[220] | p[220] &(g[219] | p[219] &(g[218] | p[218] &(g[217] | p[217] &(g[216] | p[216] &(g[215] | p[215] &(g[214] | p[214] &(g[213] | p[213] &(g[212] | p[212] &(g[211] | p[211] &(g[210] | p[210] &(g[209] | p[209] &(g[208] | p[208] &(g[207] | p[207] &(g[206] | p[206] &(g[205] | p[205] &(g[204] | p[204] &(g[203] | p[203] &(g[202] | p[202] &(g[201] | p[201] &(g[200] | p[200] &(g[199] | p[199] &(g[198] | p[198] &(g[197] | p[197] &(g[196] | p[196] &(g[195] | p[195] &(g[194] | p[194] &(g[193] | p[193] &(g[192] | p[192] &(g[191] | p[191] &(g[190] | p[190] &(g[189] | p[189] &(g[188] | p[188] &(g[187] | p[187] &(g[186] | p[186] &(g[185] | p[185] &(g[184] | p[184] &(g[183] | p[183] &(g[182] | p[182] &(g[181] | p[181] &(g[180] | p[180] &(g[179] | p[179] &(g[178] | p[178] &(g[177] | p[177] &(g[176] | p[176] &(g[175] | p[175] &(g[174] | p[174] &(g[173] | p[173] &(g[172] | p[172] &(g[171] | p[171] &(g[170] | p[170] &(g[169] | p[169] &(g[168] | p[168] &(g[167] | p[167] &(g[166] | p[166] &(g[165] | p[165] &(g[164] | p[164] &(g[163] | p[163] &(g[162] | p[162] &(g[161] | p[161] &(g[160] | p[160] &(g[159] | p[159] &(g[158] | p[158] &(g[157] | p[157] &(g[156] | p[156] &(g[155] | p[155] &(g[154] | p[154] &(g[153] | p[153] &(g[152] | p[152] &(g[151] | p[151] &(g[150] | p[150] &(g[149] | p[149] &(g[148] | p[148] &(g[147] | p[147] &(g[146] | p[146] &(g[145] | p[145] &(g[144] | p[144] &(g[143] | p[143] &(g[142] | p[142] &(g[141] | p[141] &(g[140] | p[140] &(g[139] | p[139] &(g[138] | p[138] &(g[137] | p[137] &(g[136] | p[136] &(g[135] | p[135] &(g[134] | p[134] &(g[133] | p[133] &(g[132] | p[132] &(g[131] | p[131] &(g[130] | p[130] &(g[129] | p[129] &(g[128] | p[128] &(g[127] | p[127] &(g[126] | p[126] &(g[125] | p[125] &(g[124] | p[124] &(g[123] | p[123] &(g[122] | p[122] &(g[121] | p[121] &(g[120] | p[120] &(g[119] | p[119] &(g[118] | p[118] &(g[117] | p[117] &(g[116] | p[116] &(g[115] | p[115] &(g[114] | p[114] &(g[113] | p[113] &(g[112] | p[112] &(g[111] | p[111] &(g[110] | p[110] &(g[109] | p[109] &(g[108] | p[108] &(g[107] | p[107] &(g[106] | p[106] &(g[105] | p[105] &(g[104] | p[104] &(g[103] | p[103] &(g[102] | p[102] &(g[101] | p[101] &(g[100] | p[100] &(g[99] | p[99] &(g[98] | p[98] &(g[97] | p[97] &(g[96] | p[96] &(g[95] | p[95] &(g[94] | p[94] &(g[93] | p[93] &(g[92] | p[92] &(g[91] | p[91] &(g[90] | p[90] &(g[89] | p[89] &(g[88] | p[88] &(g[87] | p[87] &(g[86] | p[86] &(g[85] | p[85] &(g[84] | p[84] &(g[83] | p[83] &(g[82] | p[82] &(g[81] | p[81] &(g[80] | p[80] &(g[79] | p[79] &(g[78] | p[78] &(g[77] | p[77] &(g[76] | p[76] &(g[75] | p[75] &(g[74] | p[74] &(g[73] | p[73] &(g[72] | p[72] &(g[71] | p[71] &(g[70] | p[70] &(g[69] | p[69] &(g[68] | p[68] &(g[67] | p[67] &(g[66] | p[66] &(g[65] | p[65] &(g[64] | p[64] &(g[63] | p[63] &(g[62] | p[62] &(g[61] | p[61] &(g[60] | p[60] &(g[59] | p[59] &(g[58] | p[58] &(g[57] | p[57] &(g[56] | p[56] &(g[55] | p[55] &(g[54] | p[54] &(g[53] | p[53] &(g[52] | p[52] &(g[51] | p[51] &(g[50] | p[50] &(g[49] | p[49] &(g[48] | p[48] &(g[47] | p[47] &(g[46] | p[46] &(g[45] | p[45] &(g[44] | p[44] &(g[43] | p[43] &(g[42] | p[42] &(g[41] | p[41] &(g[40] | p[40] &(g[39] | p[39] &(g[38] | p[38] &(g[37] | p[37] &(g[36] | p[36] &(g[35] | p[35] &(g[34] | p[34] &(g[33] | p[33] &(g[32] | p[32] &(g[31] | p[31] &(g[30] | p[30] &(g[29] | p[29] &(g[28] | p[28] &(g[27] | p[27] &(g[26] | p[26] &(g[25] | p[25] &(g[24] | p[24] &(g[23] | p[23] &(g[22] | p[22] &(g[21] | p[21] &(g[20] | p[20] &(g[19] | p[19] &(g[18] | p[18] &(g[17] | p[17] &(g[16] | p[16] &(g[15] | p[15] &(g[14] | p[14] &(g[13] | p[13] &(g[12] | p[12] &(g[11] | p[11] &(g[10] | p[10] &(g[9] | p[9] &(g[8] | p[8] &(g[7] | p[7] &(g[6] | p[6] &(g[5] | p[5] &(g[4] | p[4] &(g[3] | p[3] &(g[2] | p[2] &(g[1] | p[1] &(g[0] | carry_in[0]&p[0]))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


end
endmodule